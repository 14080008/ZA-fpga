module rom (input [16:0] address, output reg [7:0] data, output [16:0] last_address);
  assign last_address = 74161;
  always @ (*) begin
    case(address)
      17'd0: data = 8'h00;
      17'd1: data = 8'h01;
      17'd2: data = 8'h00;
      17'd3: data = 8'h02;
      17'd4: data = 8'h04;
      17'd5: data = 8'h05;
      17'd6: data = 8'h04;
      17'd7: data = 8'h05;
      17'd8: data = 8'h06;
      17'd9: data = 8'h06;
      17'd10: data = 8'h06;
      17'd11: data = 8'h0a;
      17'd12: data = 8'h0a;
      17'd13: data = 8'h09;
      17'd14: data = 8'h06;
      17'd15: data = 8'h0a;
      17'd16: data = 8'h0c;
      17'd17: data = 8'h06;
      17'd18: data = 8'h09;
      17'd19: data = 8'h09;
      17'd20: data = 8'h09;
      17'd21: data = 8'h05;
      17'd22: data = 8'h01;
      17'd23: data = 8'h02;
      17'd24: data = 8'h06;
      17'd25: data = 8'h04;
      17'd26: data = 8'h02;
      17'd27: data = 8'h05;
      17'd28: data = 8'h06;
      17'd29: data = 8'h06;
      17'd30: data = 8'h06;
      17'd31: data = 8'h0a;
      17'd32: data = 8'h0c;
      17'd33: data = 8'h05;
      17'd34: data = 8'h04;
      17'd35: data = 8'h04;
      17'd36: data = 8'h04;
      17'd37: data = 8'h02;
      17'd38: data = 8'h01;
      17'd39: data = 8'hfe;
      17'd40: data = 8'hfe;
      17'd41: data = 8'hfc;
      17'd42: data = 8'hfa;
      17'd43: data = 8'hfc;
      17'd44: data = 8'hfa;
      17'd45: data = 8'hfa;
      17'd46: data = 8'hfa;
      17'd47: data = 8'hfc;
      17'd48: data = 8'hfa;
      17'd49: data = 8'hfa;
      17'd50: data = 8'hfa;
      17'd51: data = 8'hfa;
      17'd52: data = 8'hfc;
      17'd53: data = 8'hfa;
      17'd54: data = 8'hfa;
      17'd55: data = 8'hfa;
      17'd56: data = 8'hfa;
      17'd57: data = 8'hf9;
      17'd58: data = 8'hf6;
      17'd59: data = 8'hfc;
      17'd60: data = 8'hfa;
      17'd61: data = 8'hf5;
      17'd62: data = 8'hf5;
      17'd63: data = 8'hf6;
      17'd64: data = 8'hf6;
      17'd65: data = 8'hf5;
      17'd66: data = 8'hf9;
      17'd67: data = 8'hfa;
      17'd68: data = 8'hfc;
      17'd69: data = 8'hfa;
      17'd70: data = 8'hfc;
      17'd71: data = 8'h00;
      17'd72: data = 8'h01;
      17'd73: data = 8'h00;
      17'd74: data = 8'h02;
      17'd75: data = 8'h04;
      17'd76: data = 8'h05;
      17'd77: data = 8'h06;
      17'd78: data = 8'h04;
      17'd79: data = 8'h02;
      17'd80: data = 8'h05;
      17'd81: data = 8'h04;
      17'd82: data = 8'h02;
      17'd83: data = 8'h02;
      17'd84: data = 8'h02;
      17'd85: data = 8'h04;
      17'd86: data = 8'h05;
      17'd87: data = 8'h05;
      17'd88: data = 8'h05;
      17'd89: data = 8'h05;
      17'd90: data = 8'h06;
      17'd91: data = 8'h09;
      17'd92: data = 8'h0c;
      17'd93: data = 8'h0c;
      17'd94: data = 8'h0a;
      17'd95: data = 8'h0a;
      17'd96: data = 8'h0c;
      17'd97: data = 8'h09;
      17'd98: data = 8'h06;
      17'd99: data = 8'h05;
      17'd100: data = 8'h02;
      17'd101: data = 8'h02;
      17'd102: data = 8'h01;
      17'd103: data = 8'h00;
      17'd104: data = 8'hfe;
      17'd105: data = 8'h00;
      17'd106: data = 8'h01;
      17'd107: data = 8'h01;
      17'd108: data = 8'h01;
      17'd109: data = 8'h00;
      17'd110: data = 8'h00;
      17'd111: data = 8'h00;
      17'd112: data = 8'h00;
      17'd113: data = 8'h00;
      17'd114: data = 8'hfe;
      17'd115: data = 8'hfe;
      17'd116: data = 8'hfe;
      17'd117: data = 8'h01;
      17'd118: data = 8'h02;
      17'd119: data = 8'h00;
      17'd120: data = 8'h00;
      17'd121: data = 8'hfe;
      17'd122: data = 8'hfe;
      17'd123: data = 8'hfe;
      17'd124: data = 8'hfc;
      17'd125: data = 8'hfd;
      17'd126: data = 8'hfd;
      17'd127: data = 8'hfc;
      17'd128: data = 8'hfc;
      17'd129: data = 8'hfa;
      17'd130: data = 8'hfa;
      17'd131: data = 8'hf9;
      17'd132: data = 8'hf9;
      17'd133: data = 8'hf9;
      17'd134: data = 8'hf6;
      17'd135: data = 8'hf5;
      17'd136: data = 8'hf6;
      17'd137: data = 8'hf6;
      17'd138: data = 8'hf9;
      17'd139: data = 8'hf9;
      17'd140: data = 8'hf9;
      17'd141: data = 8'hf9;
      17'd142: data = 8'hf6;
      17'd143: data = 8'hf6;
      17'd144: data = 8'hf5;
      17'd145: data = 8'hf5;
      17'd146: data = 8'hf2;
      17'd147: data = 8'hf1;
      17'd148: data = 8'hf2;
      17'd149: data = 8'hf1;
      17'd150: data = 8'hf2;
      17'd151: data = 8'hf2;
      17'd152: data = 8'hf4;
      17'd153: data = 8'hf4;
      17'd154: data = 8'hf6;
      17'd155: data = 8'hf4;
      17'd156: data = 8'hf5;
      17'd157: data = 8'hf2;
      17'd158: data = 8'hf1;
      17'd159: data = 8'hf4;
      17'd160: data = 8'hf2;
      17'd161: data = 8'hf1;
      17'd162: data = 8'hf2;
      17'd163: data = 8'hf4;
      17'd164: data = 8'hf4;
      17'd165: data = 8'hf4;
      17'd166: data = 8'hf2;
      17'd167: data = 8'hf2;
      17'd168: data = 8'hf4;
      17'd169: data = 8'hf5;
      17'd170: data = 8'hf5;
      17'd171: data = 8'hf6;
      17'd172: data = 8'hf9;
      17'd173: data = 8'hf6;
      17'd174: data = 8'hf6;
      17'd175: data = 8'hf9;
      17'd176: data = 8'hf9;
      17'd177: data = 8'hf6;
      17'd178: data = 8'hf6;
      17'd179: data = 8'hf9;
      17'd180: data = 8'hf9;
      17'd181: data = 8'hfa;
      17'd182: data = 8'hfd;
      17'd183: data = 8'h00;
      17'd184: data = 8'h02;
      17'd185: data = 8'h01;
      17'd186: data = 8'h04;
      17'd187: data = 8'h05;
      17'd188: data = 8'h02;
      17'd189: data = 8'h02;
      17'd190: data = 8'h02;
      17'd191: data = 8'h0a;
      17'd192: data = 8'h06;
      17'd193: data = 8'h00;
      17'd194: data = 8'h05;
      17'd195: data = 8'h0a;
      17'd196: data = 8'h09;
      17'd197: data = 8'h0c;
      17'd198: data = 8'h0c;
      17'd199: data = 8'h0c;
      17'd200: data = 8'h0e;
      17'd201: data = 8'h0d;
      17'd202: data = 8'h0d;
      17'd203: data = 8'h0e;
      17'd204: data = 8'h0d;
      17'd205: data = 8'h0d;
      17'd206: data = 8'h0c;
      17'd207: data = 8'h0c;
      17'd208: data = 8'h0a;
      17'd209: data = 8'h09;
      17'd210: data = 8'h0e;
      17'd211: data = 8'h0d;
      17'd212: data = 8'h0c;
      17'd213: data = 8'h0c;
      17'd214: data = 8'h0d;
      17'd215: data = 8'h11;
      17'd216: data = 8'h0e;
      17'd217: data = 8'h0a;
      17'd218: data = 8'h0c;
      17'd219: data = 8'h0a;
      17'd220: data = 8'h0a;
      17'd221: data = 8'h09;
      17'd222: data = 8'h05;
      17'd223: data = 8'h05;
      17'd224: data = 8'h09;
      17'd225: data = 8'h09;
      17'd226: data = 8'h06;
      17'd227: data = 8'h04;
      17'd228: data = 8'h02;
      17'd229: data = 8'h04;
      17'd230: data = 8'h04;
      17'd231: data = 8'h05;
      17'd232: data = 8'h04;
      17'd233: data = 8'h05;
      17'd234: data = 8'h06;
      17'd235: data = 8'h04;
      17'd236: data = 8'h05;
      17'd237: data = 8'h06;
      17'd238: data = 8'h06;
      17'd239: data = 8'h05;
      17'd240: data = 8'h04;
      17'd241: data = 8'h05;
      17'd242: data = 8'h05;
      17'd243: data = 8'h02;
      17'd244: data = 8'h05;
      17'd245: data = 8'h09;
      17'd246: data = 8'h05;
      17'd247: data = 8'h04;
      17'd248: data = 8'h06;
      17'd249: data = 8'h04;
      17'd250: data = 8'h00;
      17'd251: data = 8'hfe;
      17'd252: data = 8'h00;
      17'd253: data = 8'h04;
      17'd254: data = 8'h01;
      17'd255: data = 8'hfe;
      17'd256: data = 8'h02;
      17'd257: data = 8'h04;
      17'd258: data = 8'h04;
      17'd259: data = 8'h09;
      17'd260: data = 8'h09;
      17'd261: data = 8'h04;
      17'd262: data = 8'h01;
      17'd263: data = 8'h01;
      17'd264: data = 8'h02;
      17'd265: data = 8'h04;
      17'd266: data = 8'h00;
      17'd267: data = 8'hfd;
      17'd268: data = 8'hfc;
      17'd269: data = 8'hf9;
      17'd270: data = 8'hf6;
      17'd271: data = 8'hf6;
      17'd272: data = 8'hf5;
      17'd273: data = 8'hf4;
      17'd274: data = 8'hf4;
      17'd275: data = 8'hf4;
      17'd276: data = 8'hf5;
      17'd277: data = 8'hf4;
      17'd278: data = 8'hf5;
      17'd279: data = 8'hf6;
      17'd280: data = 8'hf5;
      17'd281: data = 8'hf6;
      17'd282: data = 8'hf6;
      17'd283: data = 8'hf6;
      17'd284: data = 8'hf4;
      17'd285: data = 8'hf1;
      17'd286: data = 8'hf2;
      17'd287: data = 8'hf2;
      17'd288: data = 8'hf1;
      17'd289: data = 8'hf1;
      17'd290: data = 8'hef;
      17'd291: data = 8'hf1;
      17'd292: data = 8'hf1;
      17'd293: data = 8'hf1;
      17'd294: data = 8'hf4;
      17'd295: data = 8'hf4;
      17'd296: data = 8'hf9;
      17'd297: data = 8'hf9;
      17'd298: data = 8'hf5;
      17'd299: data = 8'hf9;
      17'd300: data = 8'hfd;
      17'd301: data = 8'h00;
      17'd302: data = 8'hfe;
      17'd303: data = 8'h00;
      17'd304: data = 8'h02;
      17'd305: data = 8'h02;
      17'd306: data = 8'h01;
      17'd307: data = 8'h01;
      17'd308: data = 8'h01;
      17'd309: data = 8'h01;
      17'd310: data = 8'h01;
      17'd311: data = 8'h00;
      17'd312: data = 8'h00;
      17'd313: data = 8'h01;
      17'd314: data = 8'h04;
      17'd315: data = 8'h02;
      17'd316: data = 8'h02;
      17'd317: data = 8'h05;
      17'd318: data = 8'h06;
      17'd319: data = 8'h05;
      17'd320: data = 8'h05;
      17'd321: data = 8'h06;
      17'd322: data = 8'h05;
      17'd323: data = 8'h09;
      17'd324: data = 8'h06;
      17'd325: data = 8'h05;
      17'd326: data = 8'h06;
      17'd327: data = 8'h0a;
      17'd328: data = 8'h09;
      17'd329: data = 8'h04;
      17'd330: data = 8'h01;
      17'd331: data = 8'h01;
      17'd332: data = 8'h00;
      17'd333: data = 8'h00;
      17'd334: data = 8'h00;
      17'd335: data = 8'hfe;
      17'd336: data = 8'h00;
      17'd337: data = 8'h01;
      17'd338: data = 8'h02;
      17'd339: data = 8'h00;
      17'd340: data = 8'hfe;
      17'd341: data = 8'h01;
      17'd342: data = 8'h01;
      17'd343: data = 8'h00;
      17'd344: data = 8'h01;
      17'd345: data = 8'h02;
      17'd346: data = 8'h01;
      17'd347: data = 8'h01;
      17'd348: data = 8'h00;
      17'd349: data = 8'h00;
      17'd350: data = 8'hfe;
      17'd351: data = 8'hfa;
      17'd352: data = 8'hfa;
      17'd353: data = 8'hf9;
      17'd354: data = 8'hf9;
      17'd355: data = 8'hfa;
      17'd356: data = 8'hfa;
      17'd357: data = 8'hfc;
      17'd358: data = 8'hfc;
      17'd359: data = 8'hfd;
      17'd360: data = 8'hfd;
      17'd361: data = 8'hfc;
      17'd362: data = 8'hfc;
      17'd363: data = 8'hf9;
      17'd364: data = 8'hf5;
      17'd365: data = 8'hf4;
      17'd366: data = 8'hf4;
      17'd367: data = 8'hf4;
      17'd368: data = 8'hf5;
      17'd369: data = 8'hf2;
      17'd370: data = 8'hf2;
      17'd371: data = 8'hf4;
      17'd372: data = 8'hf2;
      17'd373: data = 8'hf2;
      17'd374: data = 8'hf2;
      17'd375: data = 8'hf2;
      17'd376: data = 8'hf2;
      17'd377: data = 8'hf4;
      17'd378: data = 8'hf4;
      17'd379: data = 8'hf5;
      17'd380: data = 8'hf5;
      17'd381: data = 8'hf2;
      17'd382: data = 8'hf4;
      17'd383: data = 8'hf2;
      17'd384: data = 8'hef;
      17'd385: data = 8'hed;
      17'd386: data = 8'hed;
      17'd387: data = 8'hed;
      17'd388: data = 8'hf1;
      17'd389: data = 8'hf2;
      17'd390: data = 8'hf2;
      17'd391: data = 8'hf2;
      17'd392: data = 8'hf4;
      17'd393: data = 8'hf4;
      17'd394: data = 8'hf5;
      17'd395: data = 8'hf4;
      17'd396: data = 8'hf4;
      17'd397: data = 8'hf5;
      17'd398: data = 8'hf5;
      17'd399: data = 8'hf5;
      17'd400: data = 8'hf5;
      17'd401: data = 8'hf6;
      17'd402: data = 8'hf9;
      17'd403: data = 8'hf6;
      17'd404: data = 8'hf9;
      17'd405: data = 8'hfa;
      17'd406: data = 8'hfa;
      17'd407: data = 8'hfd;
      17'd408: data = 8'hfe;
      17'd409: data = 8'hfd;
      17'd410: data = 8'hfe;
      17'd411: data = 8'h00;
      17'd412: data = 8'h01;
      17'd413: data = 8'h02;
      17'd414: data = 8'h04;
      17'd415: data = 8'h02;
      17'd416: data = 8'h05;
      17'd417: data = 8'h05;
      17'd418: data = 8'h09;
      17'd419: data = 8'h09;
      17'd420: data = 8'h05;
      17'd421: data = 8'h0c;
      17'd422: data = 8'h0e;
      17'd423: data = 8'h0d;
      17'd424: data = 8'h0e;
      17'd425: data = 8'h0e;
      17'd426: data = 8'h0d;
      17'd427: data = 8'h0c;
      17'd428: data = 8'h0a;
      17'd429: data = 8'h0a;
      17'd430: data = 8'h0c;
      17'd431: data = 8'h0a;
      17'd432: data = 8'h0c;
      17'd433: data = 8'h11;
      17'd434: data = 8'h11;
      17'd435: data = 8'h0e;
      17'd436: data = 8'h0e;
      17'd437: data = 8'h11;
      17'd438: data = 8'h0e;
      17'd439: data = 8'h0d;
      17'd440: data = 8'h0e;
      17'd441: data = 8'h11;
      17'd442: data = 8'h0c;
      17'd443: data = 8'h06;
      17'd444: data = 8'h05;
      17'd445: data = 8'h06;
      17'd446: data = 8'h06;
      17'd447: data = 8'h05;
      17'd448: data = 8'h09;
      17'd449: data = 8'h0a;
      17'd450: data = 8'h0a;
      17'd451: data = 8'h0c;
      17'd452: data = 8'h0c;
      17'd453: data = 8'h06;
      17'd454: data = 8'h0a;
      17'd455: data = 8'h0d;
      17'd456: data = 8'h0c;
      17'd457: data = 8'h09;
      17'd458: data = 8'h0c;
      17'd459: data = 8'h0a;
      17'd460: data = 8'h05;
      17'd461: data = 8'h09;
      17'd462: data = 8'h0c;
      17'd463: data = 8'h06;
      17'd464: data = 8'h01;
      17'd465: data = 8'h02;
      17'd466: data = 8'h06;
      17'd467: data = 8'h06;
      17'd468: data = 8'h04;
      17'd469: data = 8'h05;
      17'd470: data = 8'h09;
      17'd471: data = 8'h06;
      17'd472: data = 8'h06;
      17'd473: data = 8'h0d;
      17'd474: data = 8'h0d;
      17'd475: data = 8'h04;
      17'd476: data = 8'h05;
      17'd477: data = 8'h06;
      17'd478: data = 8'h06;
      17'd479: data = 8'h04;
      17'd480: data = 8'h05;
      17'd481: data = 8'h06;
      17'd482: data = 8'h02;
      17'd483: data = 8'h02;
      17'd484: data = 8'h04;
      17'd485: data = 8'h01;
      17'd486: data = 8'hfc;
      17'd487: data = 8'hf9;
      17'd488: data = 8'hf9;
      17'd489: data = 8'hfa;
      17'd490: data = 8'hf9;
      17'd491: data = 8'hf5;
      17'd492: data = 8'hf6;
      17'd493: data = 8'hf9;
      17'd494: data = 8'hf5;
      17'd495: data = 8'hf6;
      17'd496: data = 8'hf9;
      17'd497: data = 8'hf6;
      17'd498: data = 8'hf4;
      17'd499: data = 8'hf5;
      17'd500: data = 8'hf5;
      17'd501: data = 8'hf5;
      17'd502: data = 8'hf2;
      17'd503: data = 8'hf1;
      17'd504: data = 8'hf1;
      17'd505: data = 8'hef;
      17'd506: data = 8'hf1;
      17'd507: data = 8'hf1;
      17'd508: data = 8'hef;
      17'd509: data = 8'hef;
      17'd510: data = 8'hf1;
      17'd511: data = 8'hf2;
      17'd512: data = 8'hf4;
      17'd513: data = 8'hf4;
      17'd514: data = 8'hf6;
      17'd515: data = 8'hfa;
      17'd516: data = 8'hfd;
      17'd517: data = 8'h01;
      17'd518: data = 8'h01;
      17'd519: data = 8'h02;
      17'd520: data = 8'h02;
      17'd521: data = 8'h05;
      17'd522: data = 8'h05;
      17'd523: data = 8'h02;
      17'd524: data = 8'h02;
      17'd525: data = 8'h04;
      17'd526: data = 8'h01;
      17'd527: data = 8'h01;
      17'd528: data = 8'h05;
      17'd529: data = 8'h05;
      17'd530: data = 8'h04;
      17'd531: data = 8'h04;
      17'd532: data = 8'h05;
      17'd533: data = 8'h05;
      17'd534: data = 8'h05;
      17'd535: data = 8'h09;
      17'd536: data = 8'h0a;
      17'd537: data = 8'h0a;
      17'd538: data = 8'h0c;
      17'd539: data = 8'h0d;
      17'd540: data = 8'h11;
      17'd541: data = 8'h0d;
      17'd542: data = 8'h0e;
      17'd543: data = 8'h0d;
      17'd544: data = 8'h0a;
      17'd545: data = 8'h06;
      17'd546: data = 8'h04;
      17'd547: data = 8'h04;
      17'd548: data = 8'h02;
      17'd549: data = 8'h04;
      17'd550: data = 8'h04;
      17'd551: data = 8'h02;
      17'd552: data = 8'h05;
      17'd553: data = 8'h05;
      17'd554: data = 8'h02;
      17'd555: data = 8'h02;
      17'd556: data = 8'h04;
      17'd557: data = 8'h01;
      17'd558: data = 8'h00;
      17'd559: data = 8'hfe;
      17'd560: data = 8'h00;
      17'd561: data = 8'h00;
      17'd562: data = 8'h00;
      17'd563: data = 8'h02;
      17'd564: data = 8'h04;
      17'd565: data = 8'h06;
      17'd566: data = 8'h02;
      17'd567: data = 8'h00;
      17'd568: data = 8'hfd;
      17'd569: data = 8'hfc;
      17'd570: data = 8'hf6;
      17'd571: data = 8'hf4;
      17'd572: data = 8'hf5;
      17'd573: data = 8'hf5;
      17'd574: data = 8'hf6;
      17'd575: data = 8'hf6;
      17'd576: data = 8'hf9;
      17'd577: data = 8'hfa;
      17'd578: data = 8'hfa;
      17'd579: data = 8'hfc;
      17'd580: data = 8'hfa;
      17'd581: data = 8'hf5;
      17'd582: data = 8'hf6;
      17'd583: data = 8'hf6;
      17'd584: data = 8'hf2;
      17'd585: data = 8'hed;
      17'd586: data = 8'he5;
      17'd587: data = 8'hef;
      17'd588: data = 8'he9;
      17'd589: data = 8'he4;
      17'd590: data = 8'hec;
      17'd591: data = 8'hef;
      17'd592: data = 8'hec;
      17'd593: data = 8'heb;
      17'd594: data = 8'hf2;
      17'd595: data = 8'hf1;
      17'd596: data = 8'hef;
      17'd597: data = 8'hf2;
      17'd598: data = 8'hf4;
      17'd599: data = 8'hef;
      17'd600: data = 8'heb;
      17'd601: data = 8'heb;
      17'd602: data = 8'he5;
      17'd603: data = 8'he4;
      17'd604: data = 8'he9;
      17'd605: data = 8'hed;
      17'd606: data = 8'he4;
      17'd607: data = 8'he2;
      17'd608: data = 8'heb;
      17'd609: data = 8'hec;
      17'd610: data = 8'hed;
      17'd611: data = 8'hf1;
      17'd612: data = 8'hef;
      17'd613: data = 8'hef;
      17'd614: data = 8'hef;
      17'd615: data = 8'hf2;
      17'd616: data = 8'hf5;
      17'd617: data = 8'hf4;
      17'd618: data = 8'hf4;
      17'd619: data = 8'hf5;
      17'd620: data = 8'hf6;
      17'd621: data = 8'hfa;
      17'd622: data = 8'hfd;
      17'd623: data = 8'hfd;
      17'd624: data = 8'hfd;
      17'd625: data = 8'hfc;
      17'd626: data = 8'hf9;
      17'd627: data = 8'hf5;
      17'd628: data = 8'hf4;
      17'd629: data = 8'hf9;
      17'd630: data = 8'hfc;
      17'd631: data = 8'hfe;
      17'd632: data = 8'h04;
      17'd633: data = 8'h05;
      17'd634: data = 8'h05;
      17'd635: data = 8'h04;
      17'd636: data = 8'h05;
      17'd637: data = 8'h05;
      17'd638: data = 8'h06;
      17'd639: data = 8'h06;
      17'd640: data = 8'h02;
      17'd641: data = 8'h04;
      17'd642: data = 8'h0d;
      17'd643: data = 8'h11;
      17'd644: data = 8'h13;
      17'd645: data = 8'h1a;
      17'd646: data = 8'h13;
      17'd647: data = 8'h11;
      17'd648: data = 8'h0e;
      17'd649: data = 8'h0a;
      17'd650: data = 8'h09;
      17'd651: data = 8'h05;
      17'd652: data = 8'h04;
      17'd653: data = 8'h02;
      17'd654: data = 8'h02;
      17'd655: data = 8'h0a;
      17'd656: data = 8'h0d;
      17'd657: data = 8'h0d;
      17'd658: data = 8'h0e;
      17'd659: data = 8'h06;
      17'd660: data = 8'hfe;
      17'd661: data = 8'hfa;
      17'd662: data = 8'hfe;
      17'd663: data = 8'h02;
      17'd664: data = 8'h0d;
      17'd665: data = 8'h1c;
      17'd666: data = 8'h24;
      17'd667: data = 8'h29;
      17'd668: data = 8'h31;
      17'd669: data = 8'h3a;
      17'd670: data = 8'h3e;
      17'd671: data = 8'h43;
      17'd672: data = 8'h3a;
      17'd673: data = 8'h34;
      17'd674: data = 8'h2f;
      17'd675: data = 8'h2b;
      17'd676: data = 8'h2b;
      17'd677: data = 8'h2d;
      17'd678: data = 8'h2f;
      17'd679: data = 8'h22;
      17'd680: data = 8'h12;
      17'd681: data = 8'h01;
      17'd682: data = 8'hf1;
      17'd683: data = 8'he5;
      17'd684: data = 8'he2;
      17'd685: data = 8'he4;
      17'd686: data = 8'he7;
      17'd687: data = 8'he7;
      17'd688: data = 8'he7;
      17'd689: data = 8'he4;
      17'd690: data = 8'heb;
      17'd691: data = 8'hf2;
      17'd692: data = 8'hf4;
      17'd693: data = 8'hf4;
      17'd694: data = 8'he2;
      17'd695: data = 8'hd3;
      17'd696: data = 8'hca;
      17'd697: data = 8'hc6;
      17'd698: data = 8'hce;
      17'd699: data = 8'hd3;
      17'd700: data = 8'hda;
      17'd701: data = 8'hdc;
      17'd702: data = 8'hda;
      17'd703: data = 8'hdc;
      17'd704: data = 8'hde;
      17'd705: data = 8'he5;
      17'd706: data = 8'hf4;
      17'd707: data = 8'hfc;
      17'd708: data = 8'h06;
      17'd709: data = 8'h0a;
      17'd710: data = 8'h0c;
      17'd711: data = 8'h15;
      17'd712: data = 8'h1e;
      17'd713: data = 8'h27;
      17'd714: data = 8'h23;
      17'd715: data = 8'h1a;
      17'd716: data = 8'h0d;
      17'd717: data = 8'hfe;
      17'd718: data = 8'hf4;
      17'd719: data = 8'hf4;
      17'd720: data = 8'hf9;
      17'd721: data = 8'hfe;
      17'd722: data = 8'h00;
      17'd723: data = 8'hfd;
      17'd724: data = 8'h00;
      17'd725: data = 8'h04;
      17'd726: data = 8'h0a;
      17'd727: data = 8'h0e;
      17'd728: data = 8'h12;
      17'd729: data = 8'h11;
      17'd730: data = 8'h0c;
      17'd731: data = 8'h06;
      17'd732: data = 8'h06;
      17'd733: data = 8'h06;
      17'd734: data = 8'h09;
      17'd735: data = 8'h06;
      17'd736: data = 8'h04;
      17'd737: data = 8'hfd;
      17'd738: data = 8'hf9;
      17'd739: data = 8'hfa;
      17'd740: data = 8'hf9;
      17'd741: data = 8'hfc;
      17'd742: data = 8'h01;
      17'd743: data = 8'h09;
      17'd744: data = 8'h12;
      17'd745: data = 8'h22;
      17'd746: data = 8'h2b;
      17'd747: data = 8'h33;
      17'd748: data = 8'h36;
      17'd749: data = 8'h2c;
      17'd750: data = 8'h22;
      17'd751: data = 8'h12;
      17'd752: data = 8'h09;
      17'd753: data = 8'h04;
      17'd754: data = 8'h00;
      17'd755: data = 8'h00;
      17'd756: data = 8'h00;
      17'd757: data = 8'h00;
      17'd758: data = 8'h02;
      17'd759: data = 8'h05;
      17'd760: data = 8'h0d;
      17'd761: data = 8'h12;
      17'd762: data = 8'h12;
      17'd763: data = 8'h11;
      17'd764: data = 8'h0a;
      17'd765: data = 8'h05;
      17'd766: data = 8'h04;
      17'd767: data = 8'h06;
      17'd768: data = 8'h0d;
      17'd769: data = 8'h0a;
      17'd770: data = 8'h01;
      17'd771: data = 8'hfd;
      17'd772: data = 8'hf6;
      17'd773: data = 8'hf1;
      17'd774: data = 8'hf1;
      17'd775: data = 8'hf5;
      17'd776: data = 8'hfc;
      17'd777: data = 8'hfc;
      17'd778: data = 8'hfe;
      17'd779: data = 8'h01;
      17'd780: data = 8'h0c;
      17'd781: data = 8'h15;
      17'd782: data = 8'h15;
      17'd783: data = 8'h0e;
      17'd784: data = 8'h04;
      17'd785: data = 8'hf9;
      17'd786: data = 8'he9;
      17'd787: data = 8'he4;
      17'd788: data = 8'hde;
      17'd789: data = 8'hd8;
      17'd790: data = 8'hd5;
      17'd791: data = 8'hce;
      17'd792: data = 8'hca;
      17'd793: data = 8'hc9;
      17'd794: data = 8'hcb;
      17'd795: data = 8'hd1;
      17'd796: data = 8'hd6;
      17'd797: data = 8'hdc;
      17'd798: data = 8'hde;
      17'd799: data = 8'hde;
      17'd800: data = 8'he4;
      17'd801: data = 8'he7;
      17'd802: data = 8'hed;
      17'd803: data = 8'hf1;
      17'd804: data = 8'hec;
      17'd805: data = 8'he7;
      17'd806: data = 8'he3;
      17'd807: data = 8'he4;
      17'd808: data = 8'he5;
      17'd809: data = 8'heb;
      17'd810: data = 8'hf1;
      17'd811: data = 8'hf1;
      17'd812: data = 8'hf5;
      17'd813: data = 8'hfa;
      17'd814: data = 8'hfc;
      17'd815: data = 8'hfc;
      17'd816: data = 8'hf9;
      17'd817: data = 8'hf9;
      17'd818: data = 8'hf5;
      17'd819: data = 8'heb;
      17'd820: data = 8'he7;
      17'd821: data = 8'he7;
      17'd822: data = 8'heb;
      17'd823: data = 8'hf2;
      17'd824: data = 8'hf5;
      17'd825: data = 8'hf9;
      17'd826: data = 8'hf9;
      17'd827: data = 8'hf9;
      17'd828: data = 8'hfd;
      17'd829: data = 8'h02;
      17'd830: data = 8'h05;
      17'd831: data = 8'h02;
      17'd832: data = 8'h00;
      17'd833: data = 8'h02;
      17'd834: data = 8'h04;
      17'd835: data = 8'h0a;
      17'd836: data = 8'h19;
      17'd837: data = 8'h23;
      17'd838: data = 8'h1a;
      17'd839: data = 8'h15;
      17'd840: data = 8'h19;
      17'd841: data = 8'h15;
      17'd842: data = 8'h19;
      17'd843: data = 8'h1a;
      17'd844: data = 8'h1f;
      17'd845: data = 8'h16;
      17'd846: data = 8'h11;
      17'd847: data = 8'h0d;
      17'd848: data = 8'h00;
      17'd849: data = 8'h0c;
      17'd850: data = 8'hfc;
      17'd851: data = 8'h02;
      17'd852: data = 8'hf4;
      17'd853: data = 8'hf6;
      17'd854: data = 8'hec;
      17'd855: data = 8'heb;
      17'd856: data = 8'h04;
      17'd857: data = 8'h0a;
      17'd858: data = 8'h01;
      17'd859: data = 8'h09;
      17'd860: data = 8'h04;
      17'd861: data = 8'he4;
      17'd862: data = 8'hf5;
      17'd863: data = 8'h04;
      17'd864: data = 8'h12;
      17'd865: data = 8'h24;
      17'd866: data = 8'h2c;
      17'd867: data = 8'h13;
      17'd868: data = 8'hf2;
      17'd869: data = 8'hec;
      17'd870: data = 8'hd8;
      17'd871: data = 8'hd5;
      17'd872: data = 8'hd6;
      17'd873: data = 8'he9;
      17'd874: data = 8'hda;
      17'd875: data = 8'hed;
      17'd876: data = 8'h02;
      17'd877: data = 8'h00;
      17'd878: data = 8'h1b;
      17'd879: data = 8'h3a;
      17'd880: data = 8'h4a;
      17'd881: data = 8'h5a;
      17'd882: data = 8'h6c;
      17'd883: data = 8'h6a;
      17'd884: data = 8'h67;
      17'd885: data = 8'h5c;
      17'd886: data = 8'h56;
      17'd887: data = 8'h35;
      17'd888: data = 8'h1f;
      17'd889: data = 8'h09;
      17'd890: data = 8'he4;
      17'd891: data = 8'hda;
      17'd892: data = 8'hd6;
      17'd893: data = 8'hca;
      17'd894: data = 8'hc9;
      17'd895: data = 8'hd2;
      17'd896: data = 8'hd1;
      17'd897: data = 8'he2;
      17'd898: data = 8'he7;
      17'd899: data = 8'hef;
      17'd900: data = 8'hec;
      17'd901: data = 8'he2;
      17'd902: data = 8'he4;
      17'd903: data = 8'he2;
      17'd904: data = 8'hd8;
      17'd905: data = 8'hd6;
      17'd906: data = 8'hd1;
      17'd907: data = 8'hcb;
      17'd908: data = 8'hd2;
      17'd909: data = 8'hcd;
      17'd910: data = 8'he2;
      17'd911: data = 8'he9;
      17'd912: data = 8'hfc;
      17'd913: data = 8'h16;
      17'd914: data = 8'h22;
      17'd915: data = 8'h2f;
      17'd916: data = 8'h36;
      17'd917: data = 8'h35;
      17'd918: data = 8'h3a;
      17'd919: data = 8'h3d;
      17'd920: data = 8'h2f;
      17'd921: data = 8'h1e;
      17'd922: data = 8'h04;
      17'd923: data = 8'hf5;
      17'd924: data = 8'he2;
      17'd925: data = 8'he3;
      17'd926: data = 8'he4;
      17'd927: data = 8'he3;
      17'd928: data = 8'he9;
      17'd929: data = 8'hf4;
      17'd930: data = 8'hfa;
      17'd931: data = 8'h01;
      17'd932: data = 8'h11;
      17'd933: data = 8'h16;
      17'd934: data = 8'h22;
      17'd935: data = 8'h23;
      17'd936: data = 8'h23;
      17'd937: data = 8'h16;
      17'd938: data = 8'h0d;
      17'd939: data = 8'h04;
      17'd940: data = 8'hfc;
      17'd941: data = 8'hfc;
      17'd942: data = 8'hfa;
      17'd943: data = 8'hfc;
      17'd944: data = 8'hfc;
      17'd945: data = 8'h05;
      17'd946: data = 8'h0e;
      17'd947: data = 8'h1f;
      17'd948: data = 8'h2b;
      17'd949: data = 8'h35;
      17'd950: data = 8'h3a;
      17'd951: data = 8'h43;
      17'd952: data = 8'h43;
      17'd953: data = 8'h42;
      17'd954: data = 8'h35;
      17'd955: data = 8'h16;
      17'd956: data = 8'h00;
      17'd957: data = 8'heb;
      17'd958: data = 8'hd6;
      17'd959: data = 8'hd5;
      17'd960: data = 8'he4;
      17'd961: data = 8'he4;
      17'd962: data = 8'he7;
      17'd963: data = 8'hf1;
      17'd964: data = 8'hf4;
      17'd965: data = 8'hf6;
      17'd966: data = 8'hfa;
      17'd967: data = 8'h0a;
      17'd968: data = 8'h0e;
      17'd969: data = 8'h0a;
      17'd970: data = 8'h09;
      17'd971: data = 8'h02;
      17'd972: data = 8'hfc;
      17'd973: data = 8'hfd;
      17'd974: data = 8'hfa;
      17'd975: data = 8'hfd;
      17'd976: data = 8'hf4;
      17'd977: data = 8'he4;
      17'd978: data = 8'hde;
      17'd979: data = 8'he3;
      17'd980: data = 8'hec;
      17'd981: data = 8'hfc;
      17'd982: data = 8'h16;
      17'd983: data = 8'h26;
      17'd984: data = 8'h2d;
      17'd985: data = 8'h2c;
      17'd986: data = 8'h2f;
      17'd987: data = 8'h24;
      17'd988: data = 8'h12;
      17'd989: data = 8'h04;
      17'd990: data = 8'hed;
      17'd991: data = 8'hdc;
      17'd992: data = 8'hd6;
      17'd993: data = 8'hd6;
      17'd994: data = 8'hdc;
      17'd995: data = 8'hed;
      17'd996: data = 8'hf6;
      17'd997: data = 8'hfe;
      17'd998: data = 8'hfa;
      17'd999: data = 8'hf1;
      17'd1000: data = 8'heb;
      17'd1001: data = 8'he5;
      17'd1002: data = 8'he9;
      17'd1003: data = 8'he4;
      17'd1004: data = 8'he0;
      17'd1005: data = 8'hda;
      17'd1006: data = 8'hd8;
      17'd1007: data = 8'hd5;
      17'd1008: data = 8'hd8;
      17'd1009: data = 8'hda;
      17'd1010: data = 8'hdc;
      17'd1011: data = 8'he2;
      17'd1012: data = 8'he4;
      17'd1013: data = 8'hf5;
      17'd1014: data = 8'h00;
      17'd1015: data = 8'h06;
      17'd1016: data = 8'h0e;
      17'd1017: data = 8'h0c;
      17'd1018: data = 8'h01;
      17'd1019: data = 8'hf6;
      17'd1020: data = 8'he5;
      17'd1021: data = 8'hdb;
      17'd1022: data = 8'hda;
      17'd1023: data = 8'hd8;
      17'd1024: data = 8'he0;
      17'd1025: data = 8'he9;
      17'd1026: data = 8'he9;
      17'd1027: data = 8'hef;
      17'd1028: data = 8'hfc;
      17'd1029: data = 8'h04;
      17'd1030: data = 8'h01;
      17'd1031: data = 8'h00;
      17'd1032: data = 8'hfe;
      17'd1033: data = 8'hf2;
      17'd1034: data = 8'heb;
      17'd1035: data = 8'hed;
      17'd1036: data = 8'heb;
      17'd1037: data = 8'hec;
      17'd1038: data = 8'hf2;
      17'd1039: data = 8'hf1;
      17'd1040: data = 8'hf6;
      17'd1041: data = 8'hf5;
      17'd1042: data = 8'hfa;
      17'd1043: data = 8'h04;
      17'd1044: data = 8'h09;
      17'd1045: data = 8'h11;
      17'd1046: data = 8'h1a;
      17'd1047: data = 8'h15;
      17'd1048: data = 8'h13;
      17'd1049: data = 8'h12;
      17'd1050: data = 8'h13;
      17'd1051: data = 8'h16;
      17'd1052: data = 8'h05;
      17'd1053: data = 8'h00;
      17'd1054: data = 8'hfc;
      17'd1055: data = 8'hf1;
      17'd1056: data = 8'h05;
      17'd1057: data = 8'h04;
      17'd1058: data = 8'h12;
      17'd1059: data = 8'h11;
      17'd1060: data = 8'h11;
      17'd1061: data = 8'h0d;
      17'd1062: data = 8'h12;
      17'd1063: data = 8'h01;
      17'd1064: data = 8'hed;
      17'd1065: data = 8'hef;
      17'd1066: data = 8'hdc;
      17'd1067: data = 8'hd5;
      17'd1068: data = 8'hcd;
      17'd1069: data = 8'he3;
      17'd1070: data = 8'he9;
      17'd1071: data = 8'hfc;
      17'd1072: data = 8'h13;
      17'd1073: data = 8'h1c;
      17'd1074: data = 8'h16;
      17'd1075: data = 8'h1b;
      17'd1076: data = 8'h24;
      17'd1077: data = 8'h24;
      17'd1078: data = 8'h36;
      17'd1079: data = 8'h2f;
      17'd1080: data = 8'h1e;
      17'd1081: data = 8'h06;
      17'd1082: data = 8'h06;
      17'd1083: data = 8'hd8;
      17'd1084: data = 8'hb0;
      17'd1085: data = 8'haa;
      17'd1086: data = 8'h97;
      17'd1087: data = 8'h80;
      17'd1088: data = 8'h90;
      17'd1089: data = 8'hd2;
      17'd1090: data = 8'hf9;
      17'd1091: data = 8'h40;
      17'd1092: data = 8'h7f;
      17'd1093: data = 8'h7f;
      17'd1094: data = 8'h7f;
      17'd1095: data = 8'h7f;
      17'd1096: data = 8'h7f;
      17'd1097: data = 8'h4d;
      17'd1098: data = 8'h1f;
      17'd1099: data = 8'h0c;
      17'd1100: data = 8'hf6;
      17'd1101: data = 8'he9;
      17'd1102: data = 8'hdc;
      17'd1103: data = 8'hde;
      17'd1104: data = 8'h01;
      17'd1105: data = 8'h06;
      17'd1106: data = 8'h05;
      17'd1107: data = 8'h13;
      17'd1108: data = 8'h24;
      17'd1109: data = 8'h1f;
      17'd1110: data = 8'h16;
      17'd1111: data = 8'h27;
      17'd1112: data = 8'h23;
      17'd1113: data = 8'h01;
      17'd1114: data = 8'he9;
      17'd1115: data = 8'hde;
      17'd1116: data = 8'hb0;
      17'd1117: data = 8'h91;
      17'd1118: data = 8'h90;
      17'd1119: data = 8'h9a;
      17'd1120: data = 8'ha3;
      17'd1121: data = 8'hc2;
      17'd1122: data = 8'hf2;
      17'd1123: data = 8'h1a;
      17'd1124: data = 8'h39;
      17'd1125: data = 8'h5a;
      17'd1126: data = 8'h60;
      17'd1127: data = 8'h4d;
      17'd1128: data = 8'h36;
      17'd1129: data = 8'h16;
      17'd1130: data = 8'hf6;
      17'd1131: data = 8'he9;
      17'd1132: data = 8'hdb;
      17'd1133: data = 8'hce;
      17'd1134: data = 8'hcb;
      17'd1135: data = 8'hd2;
      17'd1136: data = 8'hde;
      17'd1137: data = 8'he9;
      17'd1138: data = 8'h01;
      17'd1139: data = 8'h19;
      17'd1140: data = 8'h1e;
      17'd1141: data = 8'h2d;
      17'd1142: data = 8'h34;
      17'd1143: data = 8'h29;
      17'd1144: data = 8'h22;
      17'd1145: data = 8'h1a;
      17'd1146: data = 8'h0d;
      17'd1147: data = 8'hf9;
      17'd1148: data = 8'he4;
      17'd1149: data = 8'hd2;
      17'd1150: data = 8'hc2;
      17'd1151: data = 8'hc5;
      17'd1152: data = 8'hd8;
      17'd1153: data = 8'hed;
      17'd1154: data = 8'h0e;
      17'd1155: data = 8'h29;
      17'd1156: data = 8'h35;
      17'd1157: data = 8'h45;
      17'd1158: data = 8'h4d;
      17'd1159: data = 8'h46;
      17'd1160: data = 8'h3c;
      17'd1161: data = 8'h2c;
      17'd1162: data = 8'h1b;
      17'd1163: data = 8'h02;
      17'd1164: data = 8'hf2;
      17'd1165: data = 8'hf1;
      17'd1166: data = 8'heb;
      17'd1167: data = 8'he7;
      17'd1168: data = 8'hf4;
      17'd1169: data = 8'h00;
      17'd1170: data = 8'h0c;
      17'd1171: data = 8'h1a;
      17'd1172: data = 8'h27;
      17'd1173: data = 8'h2f;
      17'd1174: data = 8'h27;
      17'd1175: data = 8'h1f;
      17'd1176: data = 8'h13;
      17'd1177: data = 8'h00;
      17'd1178: data = 8'hef;
      17'd1179: data = 8'he0;
      17'd1180: data = 8'hd3;
      17'd1181: data = 8'hcd;
      17'd1182: data = 8'hcd;
      17'd1183: data = 8'hdb;
      17'd1184: data = 8'hf1;
      17'd1185: data = 8'hfe;
      17'd1186: data = 8'h0e;
      17'd1187: data = 8'h19;
      17'd1188: data = 8'h1b;
      17'd1189: data = 8'h1f;
      17'd1190: data = 8'h1c;
      17'd1191: data = 8'h1c;
      17'd1192: data = 8'h0e;
      17'd1193: data = 8'hfc;
      17'd1194: data = 8'hf2;
      17'd1195: data = 8'he5;
      17'd1196: data = 8'hdb;
      17'd1197: data = 8'he3;
      17'd1198: data = 8'hf4;
      17'd1199: data = 8'h01;
      17'd1200: data = 8'h13;
      17'd1201: data = 8'h1e;
      17'd1202: data = 8'h1f;
      17'd1203: data = 8'h1c;
      17'd1204: data = 8'h15;
      17'd1205: data = 8'h0e;
      17'd1206: data = 8'hfe;
      17'd1207: data = 8'hf4;
      17'd1208: data = 8'he4;
      17'd1209: data = 8'hd6;
      17'd1210: data = 8'hd8;
      17'd1211: data = 8'he0;
      17'd1212: data = 8'he4;
      17'd1213: data = 8'hec;
      17'd1214: data = 8'hef;
      17'd1215: data = 8'hf2;
      17'd1216: data = 8'hf4;
      17'd1217: data = 8'hf4;
      17'd1218: data = 8'hf9;
      17'd1219: data = 8'hf1;
      17'd1220: data = 8'hf2;
      17'd1221: data = 8'hf1;
      17'd1222: data = 8'he2;
      17'd1223: data = 8'hdb;
      17'd1224: data = 8'hda;
      17'd1225: data = 8'hdc;
      17'd1226: data = 8'hde;
      17'd1227: data = 8'he3;
      17'd1228: data = 8'he9;
      17'd1229: data = 8'hef;
      17'd1230: data = 8'hfc;
      17'd1231: data = 8'hfe;
      17'd1232: data = 8'h00;
      17'd1233: data = 8'h04;
      17'd1234: data = 8'hfc;
      17'd1235: data = 8'he9;
      17'd1236: data = 8'he0;
      17'd1237: data = 8'hdb;
      17'd1238: data = 8'hd3;
      17'd1239: data = 8'hd1;
      17'd1240: data = 8'hd8;
      17'd1241: data = 8'he5;
      17'd1242: data = 8'heb;
      17'd1243: data = 8'hf5;
      17'd1244: data = 8'h01;
      17'd1245: data = 8'h00;
      17'd1246: data = 8'h02;
      17'd1247: data = 8'hf9;
      17'd1248: data = 8'hf9;
      17'd1249: data = 8'hf2;
      17'd1250: data = 8'he5;
      17'd1251: data = 8'he3;
      17'd1252: data = 8'hdc;
      17'd1253: data = 8'heb;
      17'd1254: data = 8'he7;
      17'd1255: data = 8'he4;
      17'd1256: data = 8'hf9;
      17'd1257: data = 8'hfd;
      17'd1258: data = 8'hfa;
      17'd1259: data = 8'h12;
      17'd1260: data = 8'h11;
      17'd1261: data = 8'h11;
      17'd1262: data = 8'h1e;
      17'd1263: data = 8'h1b;
      17'd1264: data = 8'h2b;
      17'd1265: data = 8'h1f;
      17'd1266: data = 8'h09;
      17'd1267: data = 8'hef;
      17'd1268: data = 8'heb;
      17'd1269: data = 8'he5;
      17'd1270: data = 8'he3;
      17'd1271: data = 8'hed;
      17'd1272: data = 8'hfd;
      17'd1273: data = 8'h06;
      17'd1274: data = 8'h0d;
      17'd1275: data = 8'h26;
      17'd1276: data = 8'h19;
      17'd1277: data = 8'h19;
      17'd1278: data = 8'h0e;
      17'd1279: data = 8'h11;
      17'd1280: data = 8'h0d;
      17'd1281: data = 8'hef;
      17'd1282: data = 8'he3;
      17'd1283: data = 8'hd3;
      17'd1284: data = 8'he3;
      17'd1285: data = 8'hef;
      17'd1286: data = 8'hf5;
      17'd1287: data = 8'hfa;
      17'd1288: data = 8'h19;
      17'd1289: data = 8'h02;
      17'd1290: data = 8'h11;
      17'd1291: data = 8'h36;
      17'd1292: data = 8'h19;
      17'd1293: data = 8'h13;
      17'd1294: data = 8'h11;
      17'd1295: data = 8'h16;
      17'd1296: data = 8'h0a;
      17'd1297: data = 8'hfc;
      17'd1298: data = 8'hc5;
      17'd1299: data = 8'h97;
      17'd1300: data = 8'h81;
      17'd1301: data = 8'h80;
      17'd1302: data = 8'haa;
      17'd1303: data = 8'hf9;
      17'd1304: data = 8'h64;
      17'd1305: data = 8'h7f;
      17'd1306: data = 8'h7f;
      17'd1307: data = 8'h7f;
      17'd1308: data = 8'h3c;
      17'd1309: data = 8'h05;
      17'd1310: data = 8'h0a;
      17'd1311: data = 8'h1e;
      17'd1312: data = 8'h33;
      17'd1313: data = 8'h27;
      17'd1314: data = 8'h1c;
      17'd1315: data = 8'h13;
      17'd1316: data = 8'hf6;
      17'd1317: data = 8'h1c;
      17'd1318: data = 8'h31;
      17'd1319: data = 8'h2f;
      17'd1320: data = 8'h2c;
      17'd1321: data = 8'h06;
      17'd1322: data = 8'h02;
      17'd1323: data = 8'h09;
      17'd1324: data = 8'h02;
      17'd1325: data = 8'h23;
      17'd1326: data = 8'h2b;
      17'd1327: data = 8'h16;
      17'd1328: data = 8'hfd;
      17'd1329: data = 8'hc0;
      17'd1330: data = 8'ha6;
      17'd1331: data = 8'h9d;
      17'd1332: data = 8'ha4;
      17'd1333: data = 8'hdb;
      17'd1334: data = 8'hf9;
      17'd1335: data = 8'h01;
      17'd1336: data = 8'h12;
      17'd1337: data = 8'h12;
      17'd1338: data = 8'h1f;
      17'd1339: data = 8'h19;
      17'd1340: data = 8'h06;
      17'd1341: data = 8'h0a;
      17'd1342: data = 8'heb;
      17'd1343: data = 8'hda;
      17'd1344: data = 8'he4;
      17'd1345: data = 8'hdb;
      17'd1346: data = 8'he9;
      17'd1347: data = 8'hed;
      17'd1348: data = 8'hf1;
      17'd1349: data = 8'h0a;
      17'd1350: data = 8'h05;
      17'd1351: data = 8'h0d;
      17'd1352: data = 8'h0c;
      17'd1353: data = 8'hfc;
      17'd1354: data = 8'h0d;
      17'd1355: data = 8'h05;
      17'd1356: data = 8'h04;
      17'd1357: data = 8'h15;
      17'd1358: data = 8'hfa;
      17'd1359: data = 8'hf6;
      17'd1360: data = 8'hf1;
      17'd1361: data = 8'hd2;
      17'd1362: data = 8'hd5;
      17'd1363: data = 8'hd5;
      17'd1364: data = 8'hec;
      17'd1365: data = 8'h0e;
      17'd1366: data = 8'h16;
      17'd1367: data = 8'h27;
      17'd1368: data = 8'h24;
      17'd1369: data = 8'h11;
      17'd1370: data = 8'h1b;
      17'd1371: data = 8'h13;
      17'd1372: data = 8'h12;
      17'd1373: data = 8'h19;
      17'd1374: data = 8'h00;
      17'd1375: data = 8'hfa;
      17'd1376: data = 8'hf9;
      17'd1377: data = 8'hf4;
      17'd1378: data = 8'h0a;
      17'd1379: data = 8'h16;
      17'd1380: data = 8'h27;
      17'd1381: data = 8'h33;
      17'd1382: data = 8'h1f;
      17'd1383: data = 8'h1c;
      17'd1384: data = 8'h0c;
      17'd1385: data = 8'h01;
      17'd1386: data = 8'h16;
      17'd1387: data = 8'h0d;
      17'd1388: data = 8'h0a;
      17'd1389: data = 8'h04;
      17'd1390: data = 8'he7;
      17'd1391: data = 8'he3;
      17'd1392: data = 8'he2;
      17'd1393: data = 8'hec;
      17'd1394: data = 8'hfe;
      17'd1395: data = 8'hf9;
      17'd1396: data = 8'hfc;
      17'd1397: data = 8'hfc;
      17'd1398: data = 8'hf5;
      17'd1399: data = 8'h04;
      17'd1400: data = 8'h0a;
      17'd1401: data = 8'h0e;
      17'd1402: data = 8'h15;
      17'd1403: data = 8'h05;
      17'd1404: data = 8'hfe;
      17'd1405: data = 8'hf9;
      17'd1406: data = 8'hf2;
      17'd1407: data = 8'hfc;
      17'd1408: data = 8'h00;
      17'd1409: data = 8'h06;
      17'd1410: data = 8'h06;
      17'd1411: data = 8'hfd;
      17'd1412: data = 8'h01;
      17'd1413: data = 8'h06;
      17'd1414: data = 8'h0a;
      17'd1415: data = 8'h16;
      17'd1416: data = 8'h15;
      17'd1417: data = 8'h0e;
      17'd1418: data = 8'h06;
      17'd1419: data = 8'hfd;
      17'd1420: data = 8'hfe;
      17'd1421: data = 8'hfd;
      17'd1422: data = 8'hf9;
      17'd1423: data = 8'hfc;
      17'd1424: data = 8'hf5;
      17'd1425: data = 8'heb;
      17'd1426: data = 8'he7;
      17'd1427: data = 8'he5;
      17'd1428: data = 8'hec;
      17'd1429: data = 8'hef;
      17'd1430: data = 8'hef;
      17'd1431: data = 8'hf2;
      17'd1432: data = 8'he9;
      17'd1433: data = 8'he7;
      17'd1434: data = 8'he9;
      17'd1435: data = 8'heb;
      17'd1436: data = 8'hf1;
      17'd1437: data = 8'he9;
      17'd1438: data = 8'he3;
      17'd1439: data = 8'he4;
      17'd1440: data = 8'he0;
      17'd1441: data = 8'he5;
      17'd1442: data = 8'hf1;
      17'd1443: data = 8'hf2;
      17'd1444: data = 8'hfa;
      17'd1445: data = 8'hf4;
      17'd1446: data = 8'hf1;
      17'd1447: data = 8'hed;
      17'd1448: data = 8'he7;
      17'd1449: data = 8'hed;
      17'd1450: data = 8'hed;
      17'd1451: data = 8'hec;
      17'd1452: data = 8'hef;
      17'd1453: data = 8'he5;
      17'd1454: data = 8'he7;
      17'd1455: data = 8'he9;
      17'd1456: data = 8'he9;
      17'd1457: data = 8'hef;
      17'd1458: data = 8'he5;
      17'd1459: data = 8'heb;
      17'd1460: data = 8'hec;
      17'd1461: data = 8'he3;
      17'd1462: data = 8'hec;
      17'd1463: data = 8'he7;
      17'd1464: data = 8'he5;
      17'd1465: data = 8'he9;
      17'd1466: data = 8'he3;
      17'd1467: data = 8'hed;
      17'd1468: data = 8'hf4;
      17'd1469: data = 8'hf9;
      17'd1470: data = 8'h0a;
      17'd1471: data = 8'h05;
      17'd1472: data = 8'h09;
      17'd1473: data = 8'h09;
      17'd1474: data = 8'h00;
      17'd1475: data = 8'h0d;
      17'd1476: data = 8'h01;
      17'd1477: data = 8'h0d;
      17'd1478: data = 8'h0a;
      17'd1479: data = 8'hfc;
      17'd1480: data = 8'h12;
      17'd1481: data = 8'h00;
      17'd1482: data = 8'hfd;
      17'd1483: data = 8'h15;
      17'd1484: data = 8'h0d;
      17'd1485: data = 8'h12;
      17'd1486: data = 8'h04;
      17'd1487: data = 8'hfe;
      17'd1488: data = 8'h09;
      17'd1489: data = 8'he7;
      17'd1490: data = 8'h0d;
      17'd1491: data = 8'h16;
      17'd1492: data = 8'hec;
      17'd1493: data = 8'h16;
      17'd1494: data = 8'h0a;
      17'd1495: data = 8'h01;
      17'd1496: data = 8'h1c;
      17'd1497: data = 8'he0;
      17'd1498: data = 8'h06;
      17'd1499: data = 8'h09;
      17'd1500: data = 8'he0;
      17'd1501: data = 8'h1c;
      17'd1502: data = 8'hed;
      17'd1503: data = 8'hda;
      17'd1504: data = 8'hf6;
      17'd1505: data = 8'hda;
      17'd1506: data = 8'h27;
      17'd1507: data = 8'h36;
      17'd1508: data = 8'h27;
      17'd1509: data = 8'h68;
      17'd1510: data = 8'h34;
      17'd1511: data = 8'h1b;
      17'd1512: data = 8'hf6;
      17'd1513: data = 8'h99;
      17'd1514: data = 8'ha4;
      17'd1515: data = 8'h83;
      17'd1516: data = 8'h91;
      17'd1517: data = 8'h05;
      17'd1518: data = 8'h1a;
      17'd1519: data = 8'h39;
      17'd1520: data = 8'h65;
      17'd1521: data = 8'h53;
      17'd1522: data = 8'h4a;
      17'd1523: data = 8'h3d;
      17'd1524: data = 8'h3e;
      17'd1525: data = 8'h3a;
      17'd1526: data = 8'h27;
      17'd1527: data = 8'h26;
      17'd1528: data = 8'h1a;
      17'd1529: data = 8'h06;
      17'd1530: data = 8'h02;
      17'd1531: data = 8'h11;
      17'd1532: data = 8'h1c;
      17'd1533: data = 8'h26;
      17'd1534: data = 8'h29;
      17'd1535: data = 8'h0a;
      17'd1536: data = 8'h19;
      17'd1537: data = 8'h22;
      17'd1538: data = 8'h19;
      17'd1539: data = 8'h2f;
      17'd1540: data = 8'h2c;
      17'd1541: data = 8'h0c;
      17'd1542: data = 8'hf5;
      17'd1543: data = 8'hd2;
      17'd1544: data = 8'hb5;
      17'd1545: data = 8'ha6;
      17'd1546: data = 8'ha6;
      17'd1547: data = 8'hca;
      17'd1548: data = 8'hdc;
      17'd1549: data = 8'hf2;
      17'd1550: data = 8'h0e;
      17'd1551: data = 8'h0d;
      17'd1552: data = 8'h0a;
      17'd1553: data = 8'h19;
      17'd1554: data = 8'h02;
      17'd1555: data = 8'hf6;
      17'd1556: data = 8'hf9;
      17'd1557: data = 8'hd8;
      17'd1558: data = 8'hd5;
      17'd1559: data = 8'hd2;
      17'd1560: data = 8'hd1;
      17'd1561: data = 8'he7;
      17'd1562: data = 8'heb;
      17'd1563: data = 8'h09;
      17'd1564: data = 8'h22;
      17'd1565: data = 8'h09;
      17'd1566: data = 8'h15;
      17'd1567: data = 8'h12;
      17'd1568: data = 8'hfe;
      17'd1569: data = 8'h11;
      17'd1570: data = 8'h11;
      17'd1571: data = 8'h0d;
      17'd1572: data = 8'h09;
      17'd1573: data = 8'he9;
      17'd1574: data = 8'he7;
      17'd1575: data = 8'he2;
      17'd1576: data = 8'hd8;
      17'd1577: data = 8'hf4;
      17'd1578: data = 8'h01;
      17'd1579: data = 8'h0d;
      17'd1580: data = 8'h22;
      17'd1581: data = 8'h1b;
      17'd1582: data = 8'h1b;
      17'd1583: data = 8'h1a;
      17'd1584: data = 8'h0e;
      17'd1585: data = 8'h12;
      17'd1586: data = 8'h0d;
      17'd1587: data = 8'hfc;
      17'd1588: data = 8'hf4;
      17'd1589: data = 8'hec;
      17'd1590: data = 8'hec;
      17'd1591: data = 8'hfe;
      17'd1592: data = 8'h06;
      17'd1593: data = 8'h23;
      17'd1594: data = 8'h35;
      17'd1595: data = 8'h2c;
      17'd1596: data = 8'h33;
      17'd1597: data = 8'h2b;
      17'd1598: data = 8'h19;
      17'd1599: data = 8'h12;
      17'd1600: data = 8'h06;
      17'd1601: data = 8'h01;
      17'd1602: data = 8'hfa;
      17'd1603: data = 8'hf6;
      17'd1604: data = 8'hf6;
      17'd1605: data = 8'hf1;
      17'd1606: data = 8'hf6;
      17'd1607: data = 8'h02;
      17'd1608: data = 8'h0c;
      17'd1609: data = 8'h0e;
      17'd1610: data = 8'h12;
      17'd1611: data = 8'h15;
      17'd1612: data = 8'h06;
      17'd1613: data = 8'h01;
      17'd1614: data = 8'h01;
      17'd1615: data = 8'hf5;
      17'd1616: data = 8'hf6;
      17'd1617: data = 8'hf1;
      17'd1618: data = 8'hed;
      17'd1619: data = 8'hf2;
      17'd1620: data = 8'hed;
      17'd1621: data = 8'h02;
      17'd1622: data = 8'h13;
      17'd1623: data = 8'h1e;
      17'd1624: data = 8'h24;
      17'd1625: data = 8'h1b;
      17'd1626: data = 8'h16;
      17'd1627: data = 8'h09;
      17'd1628: data = 8'h01;
      17'd1629: data = 8'h04;
      17'd1630: data = 8'hfe;
      17'd1631: data = 8'h00;
      17'd1632: data = 8'hfe;
      17'd1633: data = 8'h01;
      17'd1634: data = 8'h09;
      17'd1635: data = 8'hfe;
      17'd1636: data = 8'h06;
      17'd1637: data = 8'h0c;
      17'd1638: data = 8'hfc;
      17'd1639: data = 8'h05;
      17'd1640: data = 8'hf9;
      17'd1641: data = 8'hed;
      17'd1642: data = 8'hef;
      17'd1643: data = 8'hdc;
      17'd1644: data = 8'he5;
      17'd1645: data = 8'hdc;
      17'd1646: data = 8'hd1;
      17'd1647: data = 8'he0;
      17'd1648: data = 8'hd5;
      17'd1649: data = 8'he0;
      17'd1650: data = 8'hf1;
      17'd1651: data = 8'he4;
      17'd1652: data = 8'hef;
      17'd1653: data = 8'heb;
      17'd1654: data = 8'he5;
      17'd1655: data = 8'hec;
      17'd1656: data = 8'hdb;
      17'd1657: data = 8'he3;
      17'd1658: data = 8'he4;
      17'd1659: data = 8'he0;
      17'd1660: data = 8'hed;
      17'd1661: data = 8'he9;
      17'd1662: data = 8'hef;
      17'd1663: data = 8'hf4;
      17'd1664: data = 8'hf1;
      17'd1665: data = 8'hfe;
      17'd1666: data = 8'hf2;
      17'd1667: data = 8'hed;
      17'd1668: data = 8'hed;
      17'd1669: data = 8'he4;
      17'd1670: data = 8'he7;
      17'd1671: data = 8'he2;
      17'd1672: data = 8'he2;
      17'd1673: data = 8'he9;
      17'd1674: data = 8'he2;
      17'd1675: data = 8'hed;
      17'd1676: data = 8'hf4;
      17'd1677: data = 8'he7;
      17'd1678: data = 8'hed;
      17'd1679: data = 8'heb;
      17'd1680: data = 8'heb;
      17'd1681: data = 8'heb;
      17'd1682: data = 8'he3;
      17'd1683: data = 8'hf9;
      17'd1684: data = 8'hf1;
      17'd1685: data = 8'hf9;
      17'd1686: data = 8'h09;
      17'd1687: data = 8'hf6;
      17'd1688: data = 8'h05;
      17'd1689: data = 8'h13;
      17'd1690: data = 8'h12;
      17'd1691: data = 8'h1c;
      17'd1692: data = 8'h15;
      17'd1693: data = 8'h04;
      17'd1694: data = 8'h0e;
      17'd1695: data = 8'h05;
      17'd1696: data = 8'h0d;
      17'd1697: data = 8'h1c;
      17'd1698: data = 8'hf6;
      17'd1699: data = 8'h19;
      17'd1700: data = 8'h0c;
      17'd1701: data = 8'hf5;
      17'd1702: data = 8'h11;
      17'd1703: data = 8'hf5;
      17'd1704: data = 8'hfa;
      17'd1705: data = 8'h04;
      17'd1706: data = 8'h09;
      17'd1707: data = 8'h13;
      17'd1708: data = 8'h0c;
      17'd1709: data = 8'hfe;
      17'd1710: data = 8'hfc;
      17'd1711: data = 8'h00;
      17'd1712: data = 8'hfd;
      17'd1713: data = 8'heb;
      17'd1714: data = 8'h04;
      17'd1715: data = 8'h0c;
      17'd1716: data = 8'hf4;
      17'd1717: data = 8'h13;
      17'd1718: data = 8'h04;
      17'd1719: data = 8'h12;
      17'd1720: data = 8'h2c;
      17'd1721: data = 8'h05;
      17'd1722: data = 8'h3e;
      17'd1723: data = 8'h1f;
      17'd1724: data = 8'hf5;
      17'd1725: data = 8'h1e;
      17'd1726: data = 8'he2;
      17'd1727: data = 8'he7;
      17'd1728: data = 8'hde;
      17'd1729: data = 8'hab;
      17'd1730: data = 8'hd8;
      17'd1731: data = 8'hcd;
      17'd1732: data = 8'hd3;
      17'd1733: data = 8'h1b;
      17'd1734: data = 8'h29;
      17'd1735: data = 8'h54;
      17'd1736: data = 8'h75;
      17'd1737: data = 8'h70;
      17'd1738: data = 8'h75;
      17'd1739: data = 8'h42;
      17'd1740: data = 8'h26;
      17'd1741: data = 8'h13;
      17'd1742: data = 8'hfd;
      17'd1743: data = 8'hf1;
      17'd1744: data = 8'hfa;
      17'd1745: data = 8'h11;
      17'd1746: data = 8'h1f;
      17'd1747: data = 8'h3c;
      17'd1748: data = 8'h56;
      17'd1749: data = 8'h4f;
      17'd1750: data = 8'h4d;
      17'd1751: data = 8'h3e;
      17'd1752: data = 8'h1f;
      17'd1753: data = 8'h1b;
      17'd1754: data = 8'he9;
      17'd1755: data = 8'hd6;
      17'd1756: data = 8'hca;
      17'd1757: data = 8'hb3;
      17'd1758: data = 8'hb5;
      17'd1759: data = 8'hb8;
      17'd1760: data = 8'hc0;
      17'd1761: data = 8'hde;
      17'd1762: data = 8'he9;
      17'd1763: data = 8'hf4;
      17'd1764: data = 8'h12;
      17'd1765: data = 8'h00;
      17'd1766: data = 8'h02;
      17'd1767: data = 8'h00;
      17'd1768: data = 8'he5;
      17'd1769: data = 8'he0;
      17'd1770: data = 8'hc4;
      17'd1771: data = 8'hb1;
      17'd1772: data = 8'hc1;
      17'd1773: data = 8'hc0;
      17'd1774: data = 8'hce;
      17'd1775: data = 8'hf6;
      17'd1776: data = 8'h06;
      17'd1777: data = 8'h22;
      17'd1778: data = 8'h2c;
      17'd1779: data = 8'h2b;
      17'd1780: data = 8'h2c;
      17'd1781: data = 8'h16;
      17'd1782: data = 8'h05;
      17'd1783: data = 8'hfe;
      17'd1784: data = 8'hec;
      17'd1785: data = 8'he4;
      17'd1786: data = 8'he5;
      17'd1787: data = 8'hf1;
      17'd1788: data = 8'hfe;
      17'd1789: data = 8'h12;
      17'd1790: data = 8'h22;
      17'd1791: data = 8'h2c;
      17'd1792: data = 8'h33;
      17'd1793: data = 8'h2b;
      17'd1794: data = 8'h24;
      17'd1795: data = 8'h1e;
      17'd1796: data = 8'h09;
      17'd1797: data = 8'hfe;
      17'd1798: data = 8'hf6;
      17'd1799: data = 8'he7;
      17'd1800: data = 8'heb;
      17'd1801: data = 8'he5;
      17'd1802: data = 8'hef;
      17'd1803: data = 8'h02;
      17'd1804: data = 8'h0a;
      17'd1805: data = 8'h1c;
      17'd1806: data = 8'h2c;
      17'd1807: data = 8'h27;
      17'd1808: data = 8'h2b;
      17'd1809: data = 8'h22;
      17'd1810: data = 8'h0c;
      17'd1811: data = 8'h00;
      17'd1812: data = 8'hef;
      17'd1813: data = 8'he0;
      17'd1814: data = 8'he5;
      17'd1815: data = 8'hef;
      17'd1816: data = 8'hf2;
      17'd1817: data = 8'h0a;
      17'd1818: data = 8'h12;
      17'd1819: data = 8'h22;
      17'd1820: data = 8'h2f;
      17'd1821: data = 8'h23;
      17'd1822: data = 8'h26;
      17'd1823: data = 8'h1a;
      17'd1824: data = 8'hf9;
      17'd1825: data = 8'hf4;
      17'd1826: data = 8'he9;
      17'd1827: data = 8'hdb;
      17'd1828: data = 8'hed;
      17'd1829: data = 8'hef;
      17'd1830: data = 8'h05;
      17'd1831: data = 8'h1a;
      17'd1832: data = 8'h19;
      17'd1833: data = 8'h2c;
      17'd1834: data = 8'h2d;
      17'd1835: data = 8'h22;
      17'd1836: data = 8'h12;
      17'd1837: data = 8'h00;
      17'd1838: data = 8'hf9;
      17'd1839: data = 8'heb;
      17'd1840: data = 8'he5;
      17'd1841: data = 8'hf9;
      17'd1842: data = 8'hf1;
      17'd1843: data = 8'hf6;
      17'd1844: data = 8'h0c;
      17'd1845: data = 8'h0d;
      17'd1846: data = 8'h22;
      17'd1847: data = 8'h19;
      17'd1848: data = 8'h12;
      17'd1849: data = 8'h1a;
      17'd1850: data = 8'hfd;
      17'd1851: data = 8'hf1;
      17'd1852: data = 8'hef;
      17'd1853: data = 8'hd5;
      17'd1854: data = 8'hd5;
      17'd1855: data = 8'hdb;
      17'd1856: data = 8'hd5;
      17'd1857: data = 8'he7;
      17'd1858: data = 8'hec;
      17'd1859: data = 8'hed;
      17'd1860: data = 8'h02;
      17'd1861: data = 8'hfe;
      17'd1862: data = 8'hf6;
      17'd1863: data = 8'hef;
      17'd1864: data = 8'hdb;
      17'd1865: data = 8'hd2;
      17'd1866: data = 8'hca;
      17'd1867: data = 8'hcb;
      17'd1868: data = 8'hd2;
      17'd1869: data = 8'hda;
      17'd1870: data = 8'he9;
      17'd1871: data = 8'hf4;
      17'd1872: data = 8'hfe;
      17'd1873: data = 8'h01;
      17'd1874: data = 8'hfc;
      17'd1875: data = 8'hfd;
      17'd1876: data = 8'hfa;
      17'd1877: data = 8'hec;
      17'd1878: data = 8'hf2;
      17'd1879: data = 8'he5;
      17'd1880: data = 8'he0;
      17'd1881: data = 8'hf4;
      17'd1882: data = 8'he4;
      17'd1883: data = 8'hf4;
      17'd1884: data = 8'hfe;
      17'd1885: data = 8'hed;
      17'd1886: data = 8'h02;
      17'd1887: data = 8'h01;
      17'd1888: data = 8'hf5;
      17'd1889: data = 8'hf6;
      17'd1890: data = 8'hed;
      17'd1891: data = 8'hde;
      17'd1892: data = 8'hdc;
      17'd1893: data = 8'he4;
      17'd1894: data = 8'hcb;
      17'd1895: data = 8'hdb;
      17'd1896: data = 8'hef;
      17'd1897: data = 8'he0;
      17'd1898: data = 8'h0c;
      17'd1899: data = 8'h13;
      17'd1900: data = 8'hfe;
      17'd1901: data = 8'h2b;
      17'd1902: data = 8'h12;
      17'd1903: data = 8'hed;
      17'd1904: data = 8'h27;
      17'd1905: data = 8'hec;
      17'd1906: data = 8'heb;
      17'd1907: data = 8'h24;
      17'd1908: data = 8'he3;
      17'd1909: data = 8'h1e;
      17'd1910: data = 8'h2d;
      17'd1911: data = 8'hfe;
      17'd1912: data = 8'h43;
      17'd1913: data = 8'h19;
      17'd1914: data = 8'hfd;
      17'd1915: data = 8'h39;
      17'd1916: data = 8'hf5;
      17'd1917: data = 8'hf1;
      17'd1918: data = 8'h1e;
      17'd1919: data = 8'hec;
      17'd1920: data = 8'hf5;
      17'd1921: data = 8'h1b;
      17'd1922: data = 8'h15;
      17'd1923: data = 8'hef;
      17'd1924: data = 8'h00;
      17'd1925: data = 8'hf5;
      17'd1926: data = 8'hcb;
      17'd1927: data = 8'h09;
      17'd1928: data = 8'he0;
      17'd1929: data = 8'h1c;
      17'd1930: data = 8'h45;
      17'd1931: data = 8'hfa;
      17'd1932: data = 8'h42;
      17'd1933: data = 8'h36;
      17'd1934: data = 8'hdc;
      17'd1935: data = 8'h0d;
      17'd1936: data = 8'he2;
      17'd1937: data = 8'hbb;
      17'd1938: data = 8'hf1;
      17'd1939: data = 8'h9f;
      17'd1940: data = 8'he0;
      17'd1941: data = 8'h04;
      17'd1942: data = 8'hce;
      17'd1943: data = 8'h43;
      17'd1944: data = 8'h39;
      17'd1945: data = 8'h35;
      17'd1946: data = 8'h4d;
      17'd1947: data = 8'h33;
      17'd1948: data = 8'h40;
      17'd1949: data = 8'h2c;
      17'd1950: data = 8'h1b;
      17'd1951: data = 8'h26;
      17'd1952: data = 8'h0e;
      17'd1953: data = 8'h0a;
      17'd1954: data = 8'h1b;
      17'd1955: data = 8'h1f;
      17'd1956: data = 8'h40;
      17'd1957: data = 8'h40;
      17'd1958: data = 8'h6e;
      17'd1959: data = 8'h67;
      17'd1960: data = 8'h43;
      17'd1961: data = 8'h54;
      17'd1962: data = 8'h1b;
      17'd1963: data = 8'h04;
      17'd1964: data = 8'h0d;
      17'd1965: data = 8'heb;
      17'd1966: data = 8'he0;
      17'd1967: data = 8'he2;
      17'd1968: data = 8'hc5;
      17'd1969: data = 8'he2;
      17'd1970: data = 8'he5;
      17'd1971: data = 8'he2;
      17'd1972: data = 8'h0c;
      17'd1973: data = 8'hfa;
      17'd1974: data = 8'hf2;
      17'd1975: data = 8'hf9;
      17'd1976: data = 8'hd8;
      17'd1977: data = 8'hcb;
      17'd1978: data = 8'hc4;
      17'd1979: data = 8'hb5;
      17'd1980: data = 8'hc5;
      17'd1981: data = 8'hc0;
      17'd1982: data = 8'hc0;
      17'd1983: data = 8'hd3;
      17'd1984: data = 8'he3;
      17'd1985: data = 8'hf5;
      17'd1986: data = 8'h02;
      17'd1987: data = 8'h1b;
      17'd1988: data = 8'h0d;
      17'd1989: data = 8'hfe;
      17'd1990: data = 8'hfe;
      17'd1991: data = 8'heb;
      17'd1992: data = 8'he5;
      17'd1993: data = 8'he9;
      17'd1994: data = 8'he7;
      17'd1995: data = 8'hfc;
      17'd1996: data = 8'h02;
      17'd1997: data = 8'h06;
      17'd1998: data = 8'h24;
      17'd1999: data = 8'h24;
      17'd2000: data = 8'h2c;
      17'd2001: data = 8'h3c;
      17'd2002: data = 8'h2b;
      17'd2003: data = 8'h24;
      17'd2004: data = 8'h1b;
      17'd2005: data = 8'h04;
      17'd2006: data = 8'h02;
      17'd2007: data = 8'h01;
      17'd2008: data = 8'h00;
      17'd2009: data = 8'h05;
      17'd2010: data = 8'h04;
      17'd2011: data = 8'h0e;
      17'd2012: data = 8'h16;
      17'd2013: data = 8'h1a;
      17'd2014: data = 8'h1e;
      17'd2015: data = 8'h1f;
      17'd2016: data = 8'h1c;
      17'd2017: data = 8'h0e;
      17'd2018: data = 8'h05;
      17'd2019: data = 8'hfd;
      17'd2020: data = 8'he7;
      17'd2021: data = 8'he7;
      17'd2022: data = 8'hed;
      17'd2023: data = 8'hed;
      17'd2024: data = 8'hfe;
      17'd2025: data = 8'h05;
      17'd2026: data = 8'h0c;
      17'd2027: data = 8'h19;
      17'd2028: data = 8'h0e;
      17'd2029: data = 8'h11;
      17'd2030: data = 8'h11;
      17'd2031: data = 8'hfa;
      17'd2032: data = 8'hfa;
      17'd2033: data = 8'hf5;
      17'd2034: data = 8'he9;
      17'd2035: data = 8'heb;
      17'd2036: data = 8'hef;
      17'd2037: data = 8'hfc;
      17'd2038: data = 8'h02;
      17'd2039: data = 8'h0d;
      17'd2040: data = 8'h12;
      17'd2041: data = 8'h16;
      17'd2042: data = 8'h1b;
      17'd2043: data = 8'h0d;
      17'd2044: data = 8'h11;
      17'd2045: data = 8'h09;
      17'd2046: data = 8'hfc;
      17'd2047: data = 8'h01;
      17'd2048: data = 8'h00;
      17'd2049: data = 8'h01;
      17'd2050: data = 8'h0d;
      17'd2051: data = 8'h0e;
      17'd2052: data = 8'h11;
      17'd2053: data = 8'h16;
      17'd2054: data = 8'h13;
      17'd2055: data = 8'h13;
      17'd2056: data = 8'h0d;
      17'd2057: data = 8'h06;
      17'd2058: data = 8'h05;
      17'd2059: data = 8'h00;
      17'd2060: data = 8'hfa;
      17'd2061: data = 8'hf2;
      17'd2062: data = 8'hf6;
      17'd2063: data = 8'hed;
      17'd2064: data = 8'he9;
      17'd2065: data = 8'hf2;
      17'd2066: data = 8'he5;
      17'd2067: data = 8'he5;
      17'd2068: data = 8'he4;
      17'd2069: data = 8'hdc;
      17'd2070: data = 8'he2;
      17'd2071: data = 8'hd3;
      17'd2072: data = 8'hd1;
      17'd2073: data = 8'hd8;
      17'd2074: data = 8'hca;
      17'd2075: data = 8'hcb;
      17'd2076: data = 8'hd2;
      17'd2077: data = 8'hce;
      17'd2078: data = 8'hd6;
      17'd2079: data = 8'hdb;
      17'd2080: data = 8'he0;
      17'd2081: data = 8'he4;
      17'd2082: data = 8'he0;
      17'd2083: data = 8'he9;
      17'd2084: data = 8'he4;
      17'd2085: data = 8'he5;
      17'd2086: data = 8'hed;
      17'd2087: data = 8'he7;
      17'd2088: data = 8'hec;
      17'd2089: data = 8'hed;
      17'd2090: data = 8'hec;
      17'd2091: data = 8'hf6;
      17'd2092: data = 8'hf5;
      17'd2093: data = 8'hf9;
      17'd2094: data = 8'h01;
      17'd2095: data = 8'hf4;
      17'd2096: data = 8'hf9;
      17'd2097: data = 8'hfc;
      17'd2098: data = 8'he9;
      17'd2099: data = 8'hf9;
      17'd2100: data = 8'hf1;
      17'd2101: data = 8'heb;
      17'd2102: data = 8'hf9;
      17'd2103: data = 8'heb;
      17'd2104: data = 8'hef;
      17'd2105: data = 8'hf5;
      17'd2106: data = 8'hec;
      17'd2107: data = 8'hef;
      17'd2108: data = 8'hf2;
      17'd2109: data = 8'he5;
      17'd2110: data = 8'hf2;
      17'd2111: data = 8'hed;
      17'd2112: data = 8'hf2;
      17'd2113: data = 8'h0e;
      17'd2114: data = 8'hed;
      17'd2115: data = 8'h0a;
      17'd2116: data = 8'h0a;
      17'd2117: data = 8'hed;
      17'd2118: data = 8'h0e;
      17'd2119: data = 8'h06;
      17'd2120: data = 8'hfe;
      17'd2121: data = 8'h11;
      17'd2122: data = 8'h01;
      17'd2123: data = 8'h09;
      17'd2124: data = 8'h19;
      17'd2125: data = 8'h0d;
      17'd2126: data = 8'h1e;
      17'd2127: data = 8'h12;
      17'd2128: data = 8'hf2;
      17'd2129: data = 8'hfd;
      17'd2130: data = 8'hf9;
      17'd2131: data = 8'h0e;
      17'd2132: data = 8'h05;
      17'd2133: data = 8'h0c;
      17'd2134: data = 8'h39;
      17'd2135: data = 8'hf2;
      17'd2136: data = 8'h09;
      17'd2137: data = 8'h34;
      17'd2138: data = 8'hce;
      17'd2139: data = 8'h09;
      17'd2140: data = 8'h19;
      17'd2141: data = 8'hef;
      17'd2142: data = 8'h47;
      17'd2143: data = 8'hf9;
      17'd2144: data = 8'hf6;
      17'd2145: data = 8'h22;
      17'd2146: data = 8'hae;
      17'd2147: data = 8'he5;
      17'd2148: data = 8'h02;
      17'd2149: data = 8'hc5;
      17'd2150: data = 8'h04;
      17'd2151: data = 8'hef;
      17'd2152: data = 8'hfa;
      17'd2153: data = 8'h19;
      17'd2154: data = 8'hef;
      17'd2155: data = 8'h1b;
      17'd2156: data = 8'h16;
      17'd2157: data = 8'h09;
      17'd2158: data = 8'h1f;
      17'd2159: data = 8'h12;
      17'd2160: data = 8'h3e;
      17'd2161: data = 8'h2c;
      17'd2162: data = 8'h2b;
      17'd2163: data = 8'h5b;
      17'd2164: data = 8'h1a;
      17'd2165: data = 8'h29;
      17'd2166: data = 8'h36;
      17'd2167: data = 8'h12;
      17'd2168: data = 8'h42;
      17'd2169: data = 8'h3a;
      17'd2170: data = 8'h2d;
      17'd2171: data = 8'h56;
      17'd2172: data = 8'h2f;
      17'd2173: data = 8'h27;
      17'd2174: data = 8'h34;
      17'd2175: data = 8'hfd;
      17'd2176: data = 8'h01;
      17'd2177: data = 8'hfe;
      17'd2178: data = 8'hed;
      17'd2179: data = 8'hfa;
      17'd2180: data = 8'hf2;
      17'd2181: data = 8'hf2;
      17'd2182: data = 8'he9;
      17'd2183: data = 8'heb;
      17'd2184: data = 8'he7;
      17'd2185: data = 8'hd6;
      17'd2186: data = 8'hdb;
      17'd2187: data = 8'hd1;
      17'd2188: data = 8'hc5;
      17'd2189: data = 8'hce;
      17'd2190: data = 8'hcd;
      17'd2191: data = 8'hcd;
      17'd2192: data = 8'hd3;
      17'd2193: data = 8'hc6;
      17'd2194: data = 8'hc5;
      17'd2195: data = 8'hd2;
      17'd2196: data = 8'hc2;
      17'd2197: data = 8'hd5;
      17'd2198: data = 8'he7;
      17'd2199: data = 8'hd5;
      17'd2200: data = 8'hec;
      17'd2201: data = 8'hf1;
      17'd2202: data = 8'he7;
      17'd2203: data = 8'hf5;
      17'd2204: data = 8'hef;
      17'd2205: data = 8'hf6;
      17'd2206: data = 8'h04;
      17'd2207: data = 8'h02;
      17'd2208: data = 8'h11;
      17'd2209: data = 8'h1c;
      17'd2210: data = 8'h1e;
      17'd2211: data = 8'h2c;
      17'd2212: data = 8'h2c;
      17'd2213: data = 8'h2f;
      17'd2214: data = 8'h29;
      17'd2215: data = 8'h23;
      17'd2216: data = 8'h2c;
      17'd2217: data = 8'h23;
      17'd2218: data = 8'h26;
      17'd2219: data = 8'h2b;
      17'd2220: data = 8'h26;
      17'd2221: data = 8'h2d;
      17'd2222: data = 8'h29;
      17'd2223: data = 8'h23;
      17'd2224: data = 8'h26;
      17'd2225: data = 8'h1a;
      17'd2226: data = 8'h15;
      17'd2227: data = 8'h1e;
      17'd2228: data = 8'h12;
      17'd2229: data = 8'h0d;
      17'd2230: data = 8'h0d;
      17'd2231: data = 8'h02;
      17'd2232: data = 8'h01;
      17'd2233: data = 8'hf9;
      17'd2234: data = 8'hf9;
      17'd2235: data = 8'hf6;
      17'd2236: data = 8'hed;
      17'd2237: data = 8'hfa;
      17'd2238: data = 8'hf9;
      17'd2239: data = 8'hf4;
      17'd2240: data = 8'hfd;
      17'd2241: data = 8'hf1;
      17'd2242: data = 8'hf1;
      17'd2243: data = 8'hf1;
      17'd2244: data = 8'he4;
      17'd2245: data = 8'hed;
      17'd2246: data = 8'hed;
      17'd2247: data = 8'heb;
      17'd2248: data = 8'hf5;
      17'd2249: data = 8'hf9;
      17'd2250: data = 8'hf6;
      17'd2251: data = 8'hfd;
      17'd2252: data = 8'hfc;
      17'd2253: data = 8'h04;
      17'd2254: data = 8'h0c;
      17'd2255: data = 8'h09;
      17'd2256: data = 8'h0e;
      17'd2257: data = 8'h0d;
      17'd2258: data = 8'h0d;
      17'd2259: data = 8'h11;
      17'd2260: data = 8'h0d;
      17'd2261: data = 8'h19;
      17'd2262: data = 8'h15;
      17'd2263: data = 8'h12;
      17'd2264: data = 8'h1e;
      17'd2265: data = 8'h1a;
      17'd2266: data = 8'h1a;
      17'd2267: data = 8'h1c;
      17'd2268: data = 8'h15;
      17'd2269: data = 8'h16;
      17'd2270: data = 8'h12;
      17'd2271: data = 8'h0a;
      17'd2272: data = 8'h0d;
      17'd2273: data = 8'h04;
      17'd2274: data = 8'hfc;
      17'd2275: data = 8'hfc;
      17'd2276: data = 8'hf6;
      17'd2277: data = 8'hf2;
      17'd2278: data = 8'hf1;
      17'd2279: data = 8'heb;
      17'd2280: data = 8'he3;
      17'd2281: data = 8'hdc;
      17'd2282: data = 8'hd6;
      17'd2283: data = 8'hd1;
      17'd2284: data = 8'hce;
      17'd2285: data = 8'hc9;
      17'd2286: data = 8'hc4;
      17'd2287: data = 8'hc1;
      17'd2288: data = 8'hc0;
      17'd2289: data = 8'hc5;
      17'd2290: data = 8'hc4;
      17'd2291: data = 8'hc6;
      17'd2292: data = 8'hcb;
      17'd2293: data = 8'hc6;
      17'd2294: data = 8'hcb;
      17'd2295: data = 8'hd1;
      17'd2296: data = 8'hd2;
      17'd2297: data = 8'hdb;
      17'd2298: data = 8'hde;
      17'd2299: data = 8'he0;
      17'd2300: data = 8'he7;
      17'd2301: data = 8'he5;
      17'd2302: data = 8'hec;
      17'd2303: data = 8'hf2;
      17'd2304: data = 8'he9;
      17'd2305: data = 8'hfa;
      17'd2306: data = 8'h00;
      17'd2307: data = 8'hf6;
      17'd2308: data = 8'h06;
      17'd2309: data = 8'h05;
      17'd2310: data = 8'h01;
      17'd2311: data = 8'h0c;
      17'd2312: data = 8'h04;
      17'd2313: data = 8'h00;
      17'd2314: data = 8'h0c;
      17'd2315: data = 8'hfe;
      17'd2316: data = 8'h00;
      17'd2317: data = 8'h05;
      17'd2318: data = 8'hf9;
      17'd2319: data = 8'hfc;
      17'd2320: data = 8'h05;
      17'd2321: data = 8'hf2;
      17'd2322: data = 8'h02;
      17'd2323: data = 8'h0d;
      17'd2324: data = 8'hfa;
      17'd2325: data = 8'h02;
      17'd2326: data = 8'h04;
      17'd2327: data = 8'hfc;
      17'd2328: data = 8'h00;
      17'd2329: data = 8'h04;
      17'd2330: data = 8'h0a;
      17'd2331: data = 8'hf9;
      17'd2332: data = 8'hf6;
      17'd2333: data = 8'h0e;
      17'd2334: data = 8'hda;
      17'd2335: data = 8'hfa;
      17'd2336: data = 8'h1f;
      17'd2337: data = 8'he5;
      17'd2338: data = 8'h00;
      17'd2339: data = 8'h1a;
      17'd2340: data = 8'he4;
      17'd2341: data = 8'h02;
      17'd2342: data = 8'h0e;
      17'd2343: data = 8'hec;
      17'd2344: data = 8'h01;
      17'd2345: data = 8'h0d;
      17'd2346: data = 8'hfc;
      17'd2347: data = 8'h1a;
      17'd2348: data = 8'h1b;
      17'd2349: data = 8'h1b;
      17'd2350: data = 8'h0d;
      17'd2351: data = 8'h33;
      17'd2352: data = 8'h23;
      17'd2353: data = 8'he7;
      17'd2354: data = 8'h1a;
      17'd2355: data = 8'he3;
      17'd2356: data = 8'hbd;
      17'd2357: data = 8'h0c;
      17'd2358: data = 8'he0;
      17'd2359: data = 8'hf6;
      17'd2360: data = 8'h3a;
      17'd2361: data = 8'hf1;
      17'd2362: data = 8'h06;
      17'd2363: data = 8'h1f;
      17'd2364: data = 8'hf9;
      17'd2365: data = 8'h1b;
      17'd2366: data = 8'h31;
      17'd2367: data = 8'h27;
      17'd2368: data = 8'h33;
      17'd2369: data = 8'h1b;
      17'd2370: data = 8'h0e;
      17'd2371: data = 8'h0a;
      17'd2372: data = 8'h0d;
      17'd2373: data = 8'h0e;
      17'd2374: data = 8'h29;
      17'd2375: data = 8'h43;
      17'd2376: data = 8'h29;
      17'd2377: data = 8'h42;
      17'd2378: data = 8'h5a;
      17'd2379: data = 8'h2d;
      17'd2380: data = 8'h3a;
      17'd2381: data = 8'h2c;
      17'd2382: data = 8'hfd;
      17'd2383: data = 8'h11;
      17'd2384: data = 8'h06;
      17'd2385: data = 8'hf5;
      17'd2386: data = 8'h16;
      17'd2387: data = 8'h0c;
      17'd2388: data = 8'h00;
      17'd2389: data = 8'h1e;
      17'd2390: data = 8'h0d;
      17'd2391: data = 8'hed;
      17'd2392: data = 8'hf6;
      17'd2393: data = 8'he7;
      17'd2394: data = 8'he0;
      17'd2395: data = 8'hf1;
      17'd2396: data = 8'he2;
      17'd2397: data = 8'hd5;
      17'd2398: data = 8'hda;
      17'd2399: data = 8'hc4;
      17'd2400: data = 8'hc2;
      17'd2401: data = 8'hdb;
      17'd2402: data = 8'hd6;
      17'd2403: data = 8'hce;
      17'd2404: data = 8'heb;
      17'd2405: data = 8'he3;
      17'd2406: data = 8'hd8;
      17'd2407: data = 8'he4;
      17'd2408: data = 8'hd6;
      17'd2409: data = 8'hc6;
      17'd2410: data = 8'hd1;
      17'd2411: data = 8'hcd;
      17'd2412: data = 8'hd1;
      17'd2413: data = 8'he5;
      17'd2414: data = 8'he9;
      17'd2415: data = 8'hfd;
      17'd2416: data = 8'h15;
      17'd2417: data = 8'h06;
      17'd2418: data = 8'h06;
      17'd2419: data = 8'h12;
      17'd2420: data = 8'h06;
      17'd2421: data = 8'h0d;
      17'd2422: data = 8'h16;
      17'd2423: data = 8'h12;
      17'd2424: data = 8'h1a;
      17'd2425: data = 8'h23;
      17'd2426: data = 8'h24;
      17'd2427: data = 8'h2f;
      17'd2428: data = 8'h34;
      17'd2429: data = 8'h2c;
      17'd2430: data = 8'h34;
      17'd2431: data = 8'h39;
      17'd2432: data = 8'h35;
      17'd2433: data = 8'h34;
      17'd2434: data = 8'h31;
      17'd2435: data = 8'h2c;
      17'd2436: data = 8'h22;
      17'd2437: data = 8'h26;
      17'd2438: data = 8'h1e;
      17'd2439: data = 8'h1b;
      17'd2440: data = 8'h1a;
      17'd2441: data = 8'h19;
      17'd2442: data = 8'h1f;
      17'd2443: data = 8'h1e;
      17'd2444: data = 8'h16;
      17'd2445: data = 8'h13;
      17'd2446: data = 8'h06;
      17'd2447: data = 8'hfa;
      17'd2448: data = 8'hf5;
      17'd2449: data = 8'hf2;
      17'd2450: data = 8'hf1;
      17'd2451: data = 8'hec;
      17'd2452: data = 8'hef;
      17'd2453: data = 8'hf6;
      17'd2454: data = 8'hf5;
      17'd2455: data = 8'hec;
      17'd2456: data = 8'he5;
      17'd2457: data = 8'he0;
      17'd2458: data = 8'hd2;
      17'd2459: data = 8'hda;
      17'd2460: data = 8'he0;
      17'd2461: data = 8'he4;
      17'd2462: data = 8'hed;
      17'd2463: data = 8'hef;
      17'd2464: data = 8'hf2;
      17'd2465: data = 8'hf6;
      17'd2466: data = 8'hf6;
      17'd2467: data = 8'hf4;
      17'd2468: data = 8'hfc;
      17'd2469: data = 8'hfd;
      17'd2470: data = 8'h00;
      17'd2471: data = 8'h04;
      17'd2472: data = 8'h05;
      17'd2473: data = 8'h0c;
      17'd2474: data = 8'h0c;
      17'd2475: data = 8'h0e;
      17'd2476: data = 8'h12;
      17'd2477: data = 8'h15;
      17'd2478: data = 8'h1b;
      17'd2479: data = 8'h1b;
      17'd2480: data = 8'h24;
      17'd2481: data = 8'h1f;
      17'd2482: data = 8'h16;
      17'd2483: data = 8'h15;
      17'd2484: data = 8'h0c;
      17'd2485: data = 8'h04;
      17'd2486: data = 8'h05;
      17'd2487: data = 8'h00;
      17'd2488: data = 8'hfd;
      17'd2489: data = 8'h01;
      17'd2490: data = 8'hfe;
      17'd2491: data = 8'hfd;
      17'd2492: data = 8'hfa;
      17'd2493: data = 8'heb;
      17'd2494: data = 8'he3;
      17'd2495: data = 8'hde;
      17'd2496: data = 8'hce;
      17'd2497: data = 8'hd1;
      17'd2498: data = 8'hc6;
      17'd2499: data = 8'hc1;
      17'd2500: data = 8'hc2;
      17'd2501: data = 8'hc1;
      17'd2502: data = 8'hc4;
      17'd2503: data = 8'hc4;
      17'd2504: data = 8'hc0;
      17'd2505: data = 8'hc2;
      17'd2506: data = 8'hc5;
      17'd2507: data = 8'hc4;
      17'd2508: data = 8'hc9;
      17'd2509: data = 8'hc9;
      17'd2510: data = 8'hc2;
      17'd2511: data = 8'hc6;
      17'd2512: data = 8'hd3;
      17'd2513: data = 8'hd3;
      17'd2514: data = 8'hd5;
      17'd2515: data = 8'he3;
      17'd2516: data = 8'hef;
      17'd2517: data = 8'hec;
      17'd2518: data = 8'hf1;
      17'd2519: data = 8'hfd;
      17'd2520: data = 8'hf5;
      17'd2521: data = 8'hf6;
      17'd2522: data = 8'h0d;
      17'd2523: data = 8'h05;
      17'd2524: data = 8'h02;
      17'd2525: data = 8'h11;
      17'd2526: data = 8'h0d;
      17'd2527: data = 8'h0e;
      17'd2528: data = 8'h16;
      17'd2529: data = 8'h1a;
      17'd2530: data = 8'h23;
      17'd2531: data = 8'h19;
      17'd2532: data = 8'h22;
      17'd2533: data = 8'h29;
      17'd2534: data = 8'h0d;
      17'd2535: data = 8'h1a;
      17'd2536: data = 8'h13;
      17'd2537: data = 8'h0c;
      17'd2538: data = 8'h16;
      17'd2539: data = 8'h1a;
      17'd2540: data = 8'h0c;
      17'd2541: data = 8'h1c;
      17'd2542: data = 8'h0d;
      17'd2543: data = 8'hfd;
      17'd2544: data = 8'h04;
      17'd2545: data = 8'h06;
      17'd2546: data = 8'heb;
      17'd2547: data = 8'hfa;
      17'd2548: data = 8'h0a;
      17'd2549: data = 8'he4;
      17'd2550: data = 8'h0c;
      17'd2551: data = 8'h04;
      17'd2552: data = 8'he3;
      17'd2553: data = 8'h01;
      17'd2554: data = 8'hfa;
      17'd2555: data = 8'he5;
      17'd2556: data = 8'hfd;
      17'd2557: data = 8'hf5;
      17'd2558: data = 8'he5;
      17'd2559: data = 8'hfc;
      17'd2560: data = 8'h00;
      17'd2561: data = 8'hf1;
      17'd2562: data = 8'h0e;
      17'd2563: data = 8'h0c;
      17'd2564: data = 8'hfd;
      17'd2565: data = 8'h1e;
      17'd2566: data = 8'h00;
      17'd2567: data = 8'hda;
      17'd2568: data = 8'hfd;
      17'd2569: data = 8'he5;
      17'd2570: data = 8'hdb;
      17'd2571: data = 8'h1a;
      17'd2572: data = 8'h16;
      17'd2573: data = 8'h1b;
      17'd2574: data = 8'h36;
      17'd2575: data = 8'h26;
      17'd2576: data = 8'h1b;
      17'd2577: data = 8'h22;
      17'd2578: data = 8'h1a;
      17'd2579: data = 8'h11;
      17'd2580: data = 8'h13;
      17'd2581: data = 8'h1b;
      17'd2582: data = 8'h11;
      17'd2583: data = 8'h24;
      17'd2584: data = 8'h36;
      17'd2585: data = 8'h1f;
      17'd2586: data = 8'h2f;
      17'd2587: data = 8'h33;
      17'd2588: data = 8'h1c;
      17'd2589: data = 8'h3a;
      17'd2590: data = 8'h2b;
      17'd2591: data = 8'h24;
      17'd2592: data = 8'h34;
      17'd2593: data = 8'h1c;
      17'd2594: data = 8'h13;
      17'd2595: data = 8'h15;
      17'd2596: data = 8'h05;
      17'd2597: data = 8'hf6;
      17'd2598: data = 8'hfd;
      17'd2599: data = 8'h0a;
      17'd2600: data = 8'h11;
      17'd2601: data = 8'h15;
      17'd2602: data = 8'h19;
      17'd2603: data = 8'h05;
      17'd2604: data = 8'h05;
      17'd2605: data = 8'hf5;
      17'd2606: data = 8'he3;
      17'd2607: data = 8'hec;
      17'd2608: data = 8'he2;
      17'd2609: data = 8'hda;
      17'd2610: data = 8'he3;
      17'd2611: data = 8'he5;
      17'd2612: data = 8'he2;
      17'd2613: data = 8'he7;
      17'd2614: data = 8'he5;
      17'd2615: data = 8'he5;
      17'd2616: data = 8'he2;
      17'd2617: data = 8'he2;
      17'd2618: data = 8'hde;
      17'd2619: data = 8'he4;
      17'd2620: data = 8'he5;
      17'd2621: data = 8'hda;
      17'd2622: data = 8'he4;
      17'd2623: data = 8'hdc;
      17'd2624: data = 8'hd5;
      17'd2625: data = 8'he4;
      17'd2626: data = 8'heb;
      17'd2627: data = 8'hf2;
      17'd2628: data = 8'h00;
      17'd2629: data = 8'hfe;
      17'd2630: data = 8'h05;
      17'd2631: data = 8'h09;
      17'd2632: data = 8'h00;
      17'd2633: data = 8'h06;
      17'd2634: data = 8'h01;
      17'd2635: data = 8'h05;
      17'd2636: data = 8'h0d;
      17'd2637: data = 8'h15;
      17'd2638: data = 8'h23;
      17'd2639: data = 8'h1f;
      17'd2640: data = 8'h26;
      17'd2641: data = 8'h2d;
      17'd2642: data = 8'h29;
      17'd2643: data = 8'h2d;
      17'd2644: data = 8'h2d;
      17'd2645: data = 8'h27;
      17'd2646: data = 8'h2d;
      17'd2647: data = 8'h27;
      17'd2648: data = 8'h29;
      17'd2649: data = 8'h2d;
      17'd2650: data = 8'h22;
      17'd2651: data = 8'h26;
      17'd2652: data = 8'h23;
      17'd2653: data = 8'h22;
      17'd2654: data = 8'h2b;
      17'd2655: data = 8'h26;
      17'd2656: data = 8'h22;
      17'd2657: data = 8'h23;
      17'd2658: data = 8'h1a;
      17'd2659: data = 8'h13;
      17'd2660: data = 8'h0d;
      17'd2661: data = 8'h09;
      17'd2662: data = 8'h04;
      17'd2663: data = 8'hfd;
      17'd2664: data = 8'h01;
      17'd2665: data = 8'hfc;
      17'd2666: data = 8'hf9;
      17'd2667: data = 8'hf4;
      17'd2668: data = 8'heb;
      17'd2669: data = 8'heb;
      17'd2670: data = 8'heb;
      17'd2671: data = 8'he3;
      17'd2672: data = 8'he2;
      17'd2673: data = 8'he9;
      17'd2674: data = 8'he2;
      17'd2675: data = 8'he3;
      17'd2676: data = 8'he7;
      17'd2677: data = 8'he2;
      17'd2678: data = 8'he0;
      17'd2679: data = 8'he2;
      17'd2680: data = 8'he0;
      17'd2681: data = 8'he3;
      17'd2682: data = 8'he7;
      17'd2683: data = 8'he7;
      17'd2684: data = 8'hef;
      17'd2685: data = 8'hf2;
      17'd2686: data = 8'hf2;
      17'd2687: data = 8'hf9;
      17'd2688: data = 8'hfc;
      17'd2689: data = 8'hfa;
      17'd2690: data = 8'h01;
      17'd2691: data = 8'h06;
      17'd2692: data = 8'h02;
      17'd2693: data = 8'h04;
      17'd2694: data = 8'h06;
      17'd2695: data = 8'h02;
      17'd2696: data = 8'h01;
      17'd2697: data = 8'h02;
      17'd2698: data = 8'h00;
      17'd2699: data = 8'h05;
      17'd2700: data = 8'h0a;
      17'd2701: data = 8'h05;
      17'd2702: data = 8'h0d;
      17'd2703: data = 8'h06;
      17'd2704: data = 8'h01;
      17'd2705: data = 8'h04;
      17'd2706: data = 8'h00;
      17'd2707: data = 8'hfa;
      17'd2708: data = 8'hf6;
      17'd2709: data = 8'hec;
      17'd2710: data = 8'heb;
      17'd2711: data = 8'heb;
      17'd2712: data = 8'he4;
      17'd2713: data = 8'he2;
      17'd2714: data = 8'he3;
      17'd2715: data = 8'hde;
      17'd2716: data = 8'hda;
      17'd2717: data = 8'hde;
      17'd2718: data = 8'hdb;
      17'd2719: data = 8'hd6;
      17'd2720: data = 8'hd6;
      17'd2721: data = 8'hd3;
      17'd2722: data = 8'hd1;
      17'd2723: data = 8'hd1;
      17'd2724: data = 8'hce;
      17'd2725: data = 8'hd2;
      17'd2726: data = 8'hd6;
      17'd2727: data = 8'hd3;
      17'd2728: data = 8'he0;
      17'd2729: data = 8'he2;
      17'd2730: data = 8'hdc;
      17'd2731: data = 8'he9;
      17'd2732: data = 8'he2;
      17'd2733: data = 8'he5;
      17'd2734: data = 8'hed;
      17'd2735: data = 8'he5;
      17'd2736: data = 8'hec;
      17'd2737: data = 8'hfd;
      17'd2738: data = 8'h00;
      17'd2739: data = 8'h06;
      17'd2740: data = 8'h01;
      17'd2741: data = 8'h02;
      17'd2742: data = 8'h01;
      17'd2743: data = 8'h15;
      17'd2744: data = 8'h39;
      17'd2745: data = 8'h16;
      17'd2746: data = 8'hf6;
      17'd2747: data = 8'h12;
      17'd2748: data = 8'h26;
      17'd2749: data = 8'h2d;
      17'd2750: data = 8'h19;
      17'd2751: data = 8'h06;
      17'd2752: data = 8'h19;
      17'd2753: data = 8'h0e;
      17'd2754: data = 8'h1b;
      17'd2755: data = 8'h24;
      17'd2756: data = 8'h1b;
      17'd2757: data = 8'h19;
      17'd2758: data = 8'h13;
      17'd2759: data = 8'h15;
      17'd2760: data = 8'h1c;
      17'd2761: data = 8'h01;
      17'd2762: data = 8'he5;
      17'd2763: data = 8'h05;
      17'd2764: data = 8'h12;
      17'd2765: data = 8'hf9;
      17'd2766: data = 8'h05;
      17'd2767: data = 8'h0c;
      17'd2768: data = 8'h0a;
      17'd2769: data = 8'h12;
      17'd2770: data = 8'heb;
      17'd2771: data = 8'hef;
      17'd2772: data = 8'hfd;
      17'd2773: data = 8'hf1;
      17'd2774: data = 8'hfe;
      17'd2775: data = 8'hf2;
      17'd2776: data = 8'hfa;
      17'd2777: data = 8'h0d;
      17'd2778: data = 8'h02;
      17'd2779: data = 8'hf5;
      17'd2780: data = 8'hfe;
      17'd2781: data = 8'h01;
      17'd2782: data = 8'heb;
      17'd2783: data = 8'hf1;
      17'd2784: data = 8'h0d;
      17'd2785: data = 8'hf6;
      17'd2786: data = 8'hfd;
      17'd2787: data = 8'h2d;
      17'd2788: data = 8'h04;
      17'd2789: data = 8'he9;
      17'd2790: data = 8'h09;
      17'd2791: data = 8'hed;
      17'd2792: data = 8'hec;
      17'd2793: data = 8'h13;
      17'd2794: data = 8'hf5;
      17'd2795: data = 8'h02;
      17'd2796: data = 8'h23;
      17'd2797: data = 8'h1f;
      17'd2798: data = 8'h27;
      17'd2799: data = 8'h13;
      17'd2800: data = 8'hfe;
      17'd2801: data = 8'h0d;
      17'd2802: data = 8'h19;
      17'd2803: data = 8'h0d;
      17'd2804: data = 8'h0d;
      17'd2805: data = 8'h1a;
      17'd2806: data = 8'h13;
      17'd2807: data = 8'h11;
      17'd2808: data = 8'h29;
      17'd2809: data = 8'h0e;
      17'd2810: data = 8'h0a;
      17'd2811: data = 8'h29;
      17'd2812: data = 8'h13;
      17'd2813: data = 8'h15;
      17'd2814: data = 8'h2c;
      17'd2815: data = 8'h1e;
      17'd2816: data = 8'h1c;
      17'd2817: data = 8'h1c;
      17'd2818: data = 8'h09;
      17'd2819: data = 8'h05;
      17'd2820: data = 8'h06;
      17'd2821: data = 8'h06;
      17'd2822: data = 8'h11;
      17'd2823: data = 8'h19;
      17'd2824: data = 8'h0a;
      17'd2825: data = 8'h0d;
      17'd2826: data = 8'h1a;
      17'd2827: data = 8'h04;
      17'd2828: data = 8'hfe;
      17'd2829: data = 8'h00;
      17'd2830: data = 8'hef;
      17'd2831: data = 8'hfc;
      17'd2832: data = 8'h02;
      17'd2833: data = 8'hf4;
      17'd2834: data = 8'hf5;
      17'd2835: data = 8'hf6;
      17'd2836: data = 8'hed;
      17'd2837: data = 8'he5;
      17'd2838: data = 8'he4;
      17'd2839: data = 8'he3;
      17'd2840: data = 8'he5;
      17'd2841: data = 8'heb;
      17'd2842: data = 8'he5;
      17'd2843: data = 8'heb;
      17'd2844: data = 8'hed;
      17'd2845: data = 8'he5;
      17'd2846: data = 8'he3;
      17'd2847: data = 8'he4;
      17'd2848: data = 8'hdc;
      17'd2849: data = 8'he5;
      17'd2850: data = 8'hec;
      17'd2851: data = 8'he3;
      17'd2852: data = 8'hf2;
      17'd2853: data = 8'hf2;
      17'd2854: data = 8'hed;
      17'd2855: data = 8'hf1;
      17'd2856: data = 8'hf4;
      17'd2857: data = 8'hf5;
      17'd2858: data = 8'hf2;
      17'd2859: data = 8'h05;
      17'd2860: data = 8'h00;
      17'd2861: data = 8'hfc;
      17'd2862: data = 8'h12;
      17'd2863: data = 8'h05;
      17'd2864: data = 8'h05;
      17'd2865: data = 8'h0c;
      17'd2866: data = 8'h05;
      17'd2867: data = 8'h13;
      17'd2868: data = 8'h15;
      17'd2869: data = 8'h0d;
      17'd2870: data = 8'h19;
      17'd2871: data = 8'h15;
      17'd2872: data = 8'h16;
      17'd2873: data = 8'h1b;
      17'd2874: data = 8'h1a;
      17'd2875: data = 8'h19;
      17'd2876: data = 8'h15;
      17'd2877: data = 8'h16;
      17'd2878: data = 8'h13;
      17'd2879: data = 8'h19;
      17'd2880: data = 8'h19;
      17'd2881: data = 8'h0e;
      17'd2882: data = 8'h0c;
      17'd2883: data = 8'h11;
      17'd2884: data = 8'h0a;
      17'd2885: data = 8'h09;
      17'd2886: data = 8'h0a;
      17'd2887: data = 8'h09;
      17'd2888: data = 8'h04;
      17'd2889: data = 8'h02;
      17'd2890: data = 8'hfe;
      17'd2891: data = 8'hf6;
      17'd2892: data = 8'hf6;
      17'd2893: data = 8'hf1;
      17'd2894: data = 8'hef;
      17'd2895: data = 8'hef;
      17'd2896: data = 8'hed;
      17'd2897: data = 8'hf5;
      17'd2898: data = 8'hf9;
      17'd2899: data = 8'hed;
      17'd2900: data = 8'hef;
      17'd2901: data = 8'hef;
      17'd2902: data = 8'hec;
      17'd2903: data = 8'heb;
      17'd2904: data = 8'hdc;
      17'd2905: data = 8'he7;
      17'd2906: data = 8'hec;
      17'd2907: data = 8'heb;
      17'd2908: data = 8'he7;
      17'd2909: data = 8'heb;
      17'd2910: data = 8'hf2;
      17'd2911: data = 8'hec;
      17'd2912: data = 8'he7;
      17'd2913: data = 8'hf1;
      17'd2914: data = 8'hef;
      17'd2915: data = 8'hef;
      17'd2916: data = 8'hfa;
      17'd2917: data = 8'he5;
      17'd2918: data = 8'he7;
      17'd2919: data = 8'hfe;
      17'd2920: data = 8'he9;
      17'd2921: data = 8'hf4;
      17'd2922: data = 8'h0a;
      17'd2923: data = 8'hdb;
      17'd2924: data = 8'he0;
      17'd2925: data = 8'h00;
      17'd2926: data = 8'hf4;
      17'd2927: data = 8'h02;
      17'd2928: data = 8'h0e;
      17'd2929: data = 8'hb1;
      17'd2930: data = 8'heb;
      17'd2931: data = 8'h40;
      17'd2932: data = 8'hca;
      17'd2933: data = 8'hc5;
      17'd2934: data = 8'h0a;
      17'd2935: data = 8'h05;
      17'd2936: data = 8'he5;
      17'd2937: data = 8'h04;
      17'd2938: data = 8'hf4;
      17'd2939: data = 8'hab;
      17'd2940: data = 8'he7;
      17'd2941: data = 8'h3d;
      17'd2942: data = 8'h2c;
      17'd2943: data = 8'hb0;
      17'd2944: data = 8'h9d;
      17'd2945: data = 8'hf5;
      17'd2946: data = 8'h46;
      17'd2947: data = 8'h4e;
      17'd2948: data = 8'ha6;
      17'd2949: data = 8'h84;
      17'd2950: data = 8'h26;
      17'd2951: data = 8'h3c;
      17'd2952: data = 8'he0;
      17'd2953: data = 8'h3a;
      17'd2954: data = 8'hde;
      17'd2955: data = 8'h8a;
      17'd2956: data = 8'h5d;
      17'd2957: data = 8'h29;
      17'd2958: data = 8'hae;
      17'd2959: data = 8'hf4;
      17'd2960: data = 8'h1c;
      17'd2961: data = 8'h00;
      17'd2962: data = 8'hfd;
      17'd2963: data = 8'he3;
      17'd2964: data = 8'h0a;
      17'd2965: data = 8'h3a;
      17'd2966: data = 8'he4;
      17'd2967: data = 8'hda;
      17'd2968: data = 8'h0a;
      17'd2969: data = 8'h05;
      17'd2970: data = 8'h00;
      17'd2971: data = 8'h1e;
      17'd2972: data = 8'hfd;
      17'd2973: data = 8'hda;
      17'd2974: data = 8'h09;
      17'd2975: data = 8'h09;
      17'd2976: data = 8'h04;
      17'd2977: data = 8'h1a;
      17'd2978: data = 8'h1a;
      17'd2979: data = 8'hd8;
      17'd2980: data = 8'hef;
      17'd2981: data = 8'h3c;
      17'd2982: data = 8'h11;
      17'd2983: data = 8'hf2;
      17'd2984: data = 8'hf2;
      17'd2985: data = 8'hfe;
      17'd2986: data = 8'h2d;
      17'd2987: data = 8'h0c;
      17'd2988: data = 8'hec;
      17'd2989: data = 8'h09;
      17'd2990: data = 8'h13;
      17'd2991: data = 8'h2b;
      17'd2992: data = 8'h19;
      17'd2993: data = 8'hdc;
      17'd2994: data = 8'h06;
      17'd2995: data = 8'h23;
      17'd2996: data = 8'h13;
      17'd2997: data = 8'h15;
      17'd2998: data = 8'h11;
      17'd2999: data = 8'hfc;
      17'd3000: data = 8'hfa;
      17'd3001: data = 8'h1e;
      17'd3002: data = 8'h1b;
      17'd3003: data = 8'h19;
      17'd3004: data = 8'h05;
      17'd3005: data = 8'hef;
      17'd3006: data = 8'hf6;
      17'd3007: data = 8'h33;
      17'd3008: data = 8'h34;
      17'd3009: data = 8'he5;
      17'd3010: data = 8'hed;
      17'd3011: data = 8'h02;
      17'd3012: data = 8'h1a;
      17'd3013: data = 8'h24;
      17'd3014: data = 8'h02;
      17'd3015: data = 8'he2;
      17'd3016: data = 8'h01;
      17'd3017: data = 8'h1b;
      17'd3018: data = 8'h01;
      17'd3019: data = 8'h0c;
      17'd3020: data = 8'h00;
      17'd3021: data = 8'hfd;
      17'd3022: data = 8'h06;
      17'd3023: data = 8'hf6;
      17'd3024: data = 8'h06;
      17'd3025: data = 8'h1b;
      17'd3026: data = 8'hfc;
      17'd3027: data = 8'h04;
      17'd3028: data = 8'h1c;
      17'd3029: data = 8'h02;
      17'd3030: data = 8'hf2;
      17'd3031: data = 8'h05;
      17'd3032: data = 8'h19;
      17'd3033: data = 8'h0d;
      17'd3034: data = 8'hf6;
      17'd3035: data = 8'hed;
      17'd3036: data = 8'h0d;
      17'd3037: data = 8'h22;
      17'd3038: data = 8'h0c;
      17'd3039: data = 8'hf6;
      17'd3040: data = 8'hf9;
      17'd3041: data = 8'h0a;
      17'd3042: data = 8'h1a;
      17'd3043: data = 8'h06;
      17'd3044: data = 8'hf6;
      17'd3045: data = 8'hfe;
      17'd3046: data = 8'h05;
      17'd3047: data = 8'h09;
      17'd3048: data = 8'h04;
      17'd3049: data = 8'h01;
      17'd3050: data = 8'h00;
      17'd3051: data = 8'h06;
      17'd3052: data = 8'h04;
      17'd3053: data = 8'h01;
      17'd3054: data = 8'h0a;
      17'd3055: data = 8'h00;
      17'd3056: data = 8'h05;
      17'd3057: data = 8'h16;
      17'd3058: data = 8'h02;
      17'd3059: data = 8'hf5;
      17'd3060: data = 8'h01;
      17'd3061: data = 8'h06;
      17'd3062: data = 8'h06;
      17'd3063: data = 8'h00;
      17'd3064: data = 8'hf5;
      17'd3065: data = 8'hf5;
      17'd3066: data = 8'h04;
      17'd3067: data = 8'h09;
      17'd3068: data = 8'hfd;
      17'd3069: data = 8'hf5;
      17'd3070: data = 8'hf6;
      17'd3071: data = 8'hf6;
      17'd3072: data = 8'h05;
      17'd3073: data = 8'hfd;
      17'd3074: data = 8'hf2;
      17'd3075: data = 8'hf9;
      17'd3076: data = 8'hf4;
      17'd3077: data = 8'hfa;
      17'd3078: data = 8'hf4;
      17'd3079: data = 8'hed;
      17'd3080: data = 8'hfc;
      17'd3081: data = 8'hf1;
      17'd3082: data = 8'he7;
      17'd3083: data = 8'hfc;
      17'd3084: data = 8'h00;
      17'd3085: data = 8'he9;
      17'd3086: data = 8'hf1;
      17'd3087: data = 8'h0e;
      17'd3088: data = 8'hf6;
      17'd3089: data = 8'hd5;
      17'd3090: data = 8'hfc;
      17'd3091: data = 8'hfd;
      17'd3092: data = 8'heb;
      17'd3093: data = 8'hfc;
      17'd3094: data = 8'he3;
      17'd3095: data = 8'he3;
      17'd3096: data = 8'h0d;
      17'd3097: data = 8'hfe;
      17'd3098: data = 8'hed;
      17'd3099: data = 8'hf4;
      17'd3100: data = 8'hf1;
      17'd3101: data = 8'h00;
      17'd3102: data = 8'h0a;
      17'd3103: data = 8'hfd;
      17'd3104: data = 8'hec;
      17'd3105: data = 8'hf1;
      17'd3106: data = 8'h04;
      17'd3107: data = 8'h09;
      17'd3108: data = 8'h01;
      17'd3109: data = 8'heb;
      17'd3110: data = 8'he5;
      17'd3111: data = 8'h06;
      17'd3112: data = 8'h1a;
      17'd3113: data = 8'hfc;
      17'd3114: data = 8'hec;
      17'd3115: data = 8'hfe;
      17'd3116: data = 8'h04;
      17'd3117: data = 8'h09;
      17'd3118: data = 8'hfc;
      17'd3119: data = 8'hf6;
      17'd3120: data = 8'hfd;
      17'd3121: data = 8'hf1;
      17'd3122: data = 8'h05;
      17'd3123: data = 8'h0e;
      17'd3124: data = 8'hef;
      17'd3125: data = 8'hf9;
      17'd3126: data = 8'h12;
      17'd3127: data = 8'h0a;
      17'd3128: data = 8'hf6;
      17'd3129: data = 8'hfc;
      17'd3130: data = 8'h05;
      17'd3131: data = 8'h05;
      17'd3132: data = 8'h00;
      17'd3133: data = 8'hf4;
      17'd3134: data = 8'h09;
      17'd3135: data = 8'h11;
      17'd3136: data = 8'he5;
      17'd3137: data = 8'hf9;
      17'd3138: data = 8'h1b;
      17'd3139: data = 8'h02;
      17'd3140: data = 8'hf4;
      17'd3141: data = 8'hf6;
      17'd3142: data = 8'h0d;
      17'd3143: data = 8'hfa;
      17'd3144: data = 8'hec;
      17'd3145: data = 8'h06;
      17'd3146: data = 8'hf4;
      17'd3147: data = 8'hec;
      17'd3148: data = 8'hf6;
      17'd3149: data = 8'hfd;
      17'd3150: data = 8'h0d;
      17'd3151: data = 8'hf6;
      17'd3152: data = 8'hd3;
      17'd3153: data = 8'h05;
      17'd3154: data = 8'h0c;
      17'd3155: data = 8'he3;
      17'd3156: data = 8'hfe;
      17'd3157: data = 8'hfa;
      17'd3158: data = 8'hed;
      17'd3159: data = 8'hfc;
      17'd3160: data = 8'hec;
      17'd3161: data = 8'hf6;
      17'd3162: data = 8'h31;
      17'd3163: data = 8'hef;
      17'd3164: data = 8'hbb;
      17'd3165: data = 8'h1c;
      17'd3166: data = 8'h01;
      17'd3167: data = 8'h01;
      17'd3168: data = 8'h19;
      17'd3169: data = 8'hbc;
      17'd3170: data = 8'hed;
      17'd3171: data = 8'h31;
      17'd3172: data = 8'hfc;
      17'd3173: data = 8'hde;
      17'd3174: data = 8'hed;
      17'd3175: data = 8'hf9;
      17'd3176: data = 8'h1f;
      17'd3177: data = 8'heb;
      17'd3178: data = 8'hf4;
      17'd3179: data = 8'h23;
      17'd3180: data = 8'hda;
      17'd3181: data = 8'hf1;
      17'd3182: data = 8'h0a;
      17'd3183: data = 8'hfa;
      17'd3184: data = 8'hfd;
      17'd3185: data = 8'he0;
      17'd3186: data = 8'he9;
      17'd3187: data = 8'h11;
      17'd3188: data = 8'h12;
      17'd3189: data = 8'he7;
      17'd3190: data = 8'hcd;
      17'd3191: data = 8'h23;
      17'd3192: data = 8'h1b;
      17'd3193: data = 8'hce;
      17'd3194: data = 8'he3;
      17'd3195: data = 8'h0e;
      17'd3196: data = 8'h1c;
      17'd3197: data = 8'he7;
      17'd3198: data = 8'hce;
      17'd3199: data = 8'h13;
      17'd3200: data = 8'h12;
      17'd3201: data = 8'h00;
      17'd3202: data = 8'hf2;
      17'd3203: data = 8'he3;
      17'd3204: data = 8'h22;
      17'd3205: data = 8'h1c;
      17'd3206: data = 8'hfa;
      17'd3207: data = 8'he5;
      17'd3208: data = 8'h15;
      17'd3209: data = 8'h26;
      17'd3210: data = 8'he7;
      17'd3211: data = 8'h01;
      17'd3212: data = 8'h1c;
      17'd3213: data = 8'h04;
      17'd3214: data = 8'hf9;
      17'd3215: data = 8'h24;
      17'd3216: data = 8'h12;
      17'd3217: data = 8'hf1;
      17'd3218: data = 8'h15;
      17'd3219: data = 8'h0d;
      17'd3220: data = 8'h0a;
      17'd3221: data = 8'h19;
      17'd3222: data = 8'h02;
      17'd3223: data = 8'h02;
      17'd3224: data = 8'h0e;
      17'd3225: data = 8'h05;
      17'd3226: data = 8'h11;
      17'd3227: data = 8'h09;
      17'd3228: data = 8'hf2;
      17'd3229: data = 8'h1e;
      17'd3230: data = 8'h29;
      17'd3231: data = 8'hd3;
      17'd3232: data = 8'hf9;
      17'd3233: data = 8'h3a;
      17'd3234: data = 8'h0c;
      17'd3235: data = 8'h0a;
      17'd3236: data = 8'hf1;
      17'd3237: data = 8'hef;
      17'd3238: data = 8'h26;
      17'd3239: data = 8'h1b;
      17'd3240: data = 8'h01;
      17'd3241: data = 8'he0;
      17'd3242: data = 8'hfa;
      17'd3243: data = 8'h27;
      17'd3244: data = 8'hfc;
      17'd3245: data = 8'h01;
      17'd3246: data = 8'h15;
      17'd3247: data = 8'he9;
      17'd3248: data = 8'hf6;
      17'd3249: data = 8'h22;
      17'd3250: data = 8'h16;
      17'd3251: data = 8'hfa;
      17'd3252: data = 8'hef;
      17'd3253: data = 8'hfa;
      17'd3254: data = 8'h12;
      17'd3255: data = 8'h11;
      17'd3256: data = 8'hf4;
      17'd3257: data = 8'he7;
      17'd3258: data = 8'h09;
      17'd3259: data = 8'h04;
      17'd3260: data = 8'h02;
      17'd3261: data = 8'h06;
      17'd3262: data = 8'he3;
      17'd3263: data = 8'h11;
      17'd3264: data = 8'h0a;
      17'd3265: data = 8'h0a;
      17'd3266: data = 8'h00;
      17'd3267: data = 8'hce;
      17'd3268: data = 8'h24;
      17'd3269: data = 8'h24;
      17'd3270: data = 8'hd3;
      17'd3271: data = 8'hf1;
      17'd3272: data = 8'h11;
      17'd3273: data = 8'h16;
      17'd3274: data = 8'h01;
      17'd3275: data = 8'hc2;
      17'd3276: data = 8'h05;
      17'd3277: data = 8'h31;
      17'd3278: data = 8'hef;
      17'd3279: data = 8'hec;
      17'd3280: data = 8'hfc;
      17'd3281: data = 8'h0d;
      17'd3282: data = 8'h04;
      17'd3283: data = 8'hf1;
      17'd3284: data = 8'h09;
      17'd3285: data = 8'h02;
      17'd3286: data = 8'hf1;
      17'd3287: data = 8'hfd;
      17'd3288: data = 8'h02;
      17'd3289: data = 8'h05;
      17'd3290: data = 8'he7;
      17'd3291: data = 8'hec;
      17'd3292: data = 8'h0c;
      17'd3293: data = 8'h0e;
      17'd3294: data = 8'hf1;
      17'd3295: data = 8'hf2;
      17'd3296: data = 8'h0c;
      17'd3297: data = 8'h04;
      17'd3298: data = 8'hf1;
      17'd3299: data = 8'h09;
      17'd3300: data = 8'h06;
      17'd3301: data = 8'he4;
      17'd3302: data = 8'h0d;
      17'd3303: data = 8'hfe;
      17'd3304: data = 8'he5;
      17'd3305: data = 8'h11;
      17'd3306: data = 8'hf1;
      17'd3307: data = 8'hfa;
      17'd3308: data = 8'h1c;
      17'd3309: data = 8'hef;
      17'd3310: data = 8'hfe;
      17'd3311: data = 8'h0c;
      17'd3312: data = 8'hfa;
      17'd3313: data = 8'h04;
      17'd3314: data = 8'h04;
      17'd3315: data = 8'h13;
      17'd3316: data = 8'hf6;
      17'd3317: data = 8'he7;
      17'd3318: data = 8'h19;
      17'd3319: data = 8'h0c;
      17'd3320: data = 8'hfc;
      17'd3321: data = 8'hfa;
      17'd3322: data = 8'h02;
      17'd3323: data = 8'h1e;
      17'd3324: data = 8'hfa;
      17'd3325: data = 8'hf5;
      17'd3326: data = 8'h11;
      17'd3327: data = 8'h06;
      17'd3328: data = 8'h05;
      17'd3329: data = 8'hef;
      17'd3330: data = 8'hfd;
      17'd3331: data = 8'h0a;
      17'd3332: data = 8'h0a;
      17'd3333: data = 8'hf9;
      17'd3334: data = 8'he0;
      17'd3335: data = 8'h15;
      17'd3336: data = 8'h1b;
      17'd3337: data = 8'hf5;
      17'd3338: data = 8'hfc;
      17'd3339: data = 8'hfa;
      17'd3340: data = 8'h09;
      17'd3341: data = 8'h12;
      17'd3342: data = 8'hfc;
      17'd3343: data = 8'hfa;
      17'd3344: data = 8'hf2;
      17'd3345: data = 8'h16;
      17'd3346: data = 8'h00;
      17'd3347: data = 8'he5;
      17'd3348: data = 8'h15;
      17'd3349: data = 8'h06;
      17'd3350: data = 8'he5;
      17'd3351: data = 8'h00;
      17'd3352: data = 8'h0a;
      17'd3353: data = 8'h00;
      17'd3354: data = 8'h0e;
      17'd3355: data = 8'he2;
      17'd3356: data = 8'hf9;
      17'd3357: data = 8'h19;
      17'd3358: data = 8'hfe;
      17'd3359: data = 8'hfa;
      17'd3360: data = 8'hf4;
      17'd3361: data = 8'hfc;
      17'd3362: data = 8'h0c;
      17'd3363: data = 8'heb;
      17'd3364: data = 8'hf9;
      17'd3365: data = 8'h24;
      17'd3366: data = 8'hdb;
      17'd3367: data = 8'heb;
      17'd3368: data = 8'h1b;
      17'd3369: data = 8'hfe;
      17'd3370: data = 8'heb;
      17'd3371: data = 8'h0a;
      17'd3372: data = 8'hfe;
      17'd3373: data = 8'he9;
      17'd3374: data = 8'h12;
      17'd3375: data = 8'h0d;
      17'd3376: data = 8'he7;
      17'd3377: data = 8'he4;
      17'd3378: data = 8'h19;
      17'd3379: data = 8'h11;
      17'd3380: data = 8'heb;
      17'd3381: data = 8'hed;
      17'd3382: data = 8'h0e;
      17'd3383: data = 8'hfc;
      17'd3384: data = 8'hf5;
      17'd3385: data = 8'h1a;
      17'd3386: data = 8'he4;
      17'd3387: data = 8'hec;
      17'd3388: data = 8'h13;
      17'd3389: data = 8'hfa;
      17'd3390: data = 8'hf6;
      17'd3391: data = 8'h01;
      17'd3392: data = 8'hf4;
      17'd3393: data = 8'hed;
      17'd3394: data = 8'h0a;
      17'd3395: data = 8'h0c;
      17'd3396: data = 8'he7;
      17'd3397: data = 8'heb;
      17'd3398: data = 8'h0a;
      17'd3399: data = 8'h02;
      17'd3400: data = 8'he9;
      17'd3401: data = 8'hf6;
      17'd3402: data = 8'h12;
      17'd3403: data = 8'he7;
      17'd3404: data = 8'hf1;
      17'd3405: data = 8'h09;
      17'd3406: data = 8'hf5;
      17'd3407: data = 8'hfc;
      17'd3408: data = 8'hf1;
      17'd3409: data = 8'h00;
      17'd3410: data = 8'h00;
      17'd3411: data = 8'hfc;
      17'd3412: data = 8'hf9;
      17'd3413: data = 8'hfa;
      17'd3414: data = 8'hf2;
      17'd3415: data = 8'h16;
      17'd3416: data = 8'h09;
      17'd3417: data = 8'he2;
      17'd3418: data = 8'hef;
      17'd3419: data = 8'h0d;
      17'd3420: data = 8'h2d;
      17'd3421: data = 8'hd3;
      17'd3422: data = 8'h00;
      17'd3423: data = 8'h2b;
      17'd3424: data = 8'he4;
      17'd3425: data = 8'h0e;
      17'd3426: data = 8'h06;
      17'd3427: data = 8'hfa;
      17'd3428: data = 8'h15;
      17'd3429: data = 8'hfd;
      17'd3430: data = 8'hf6;
      17'd3431: data = 8'h16;
      17'd3432: data = 8'h09;
      17'd3433: data = 8'h02;
      17'd3434: data = 8'hf9;
      17'd3435: data = 8'h02;
      17'd3436: data = 8'h1e;
      17'd3437: data = 8'h11;
      17'd3438: data = 8'he3;
      17'd3439: data = 8'hfa;
      17'd3440: data = 8'h33;
      17'd3441: data = 8'h04;
      17'd3442: data = 8'he3;
      17'd3443: data = 8'h16;
      17'd3444: data = 8'hf5;
      17'd3445: data = 8'h00;
      17'd3446: data = 8'h2f;
      17'd3447: data = 8'hdc;
      17'd3448: data = 8'hed;
      17'd3449: data = 8'h29;
      17'd3450: data = 8'hfe;
      17'd3451: data = 8'hf6;
      17'd3452: data = 8'hf9;
      17'd3453: data = 8'h13;
      17'd3454: data = 8'h0c;
      17'd3455: data = 8'he5;
      17'd3456: data = 8'h19;
      17'd3457: data = 8'hf9;
      17'd3458: data = 8'h00;
      17'd3459: data = 8'h00;
      17'd3460: data = 8'hf2;
      17'd3461: data = 8'h29;
      17'd3462: data = 8'he2;
      17'd3463: data = 8'hed;
      17'd3464: data = 8'h0e;
      17'd3465: data = 8'h04;
      17'd3466: data = 8'h19;
      17'd3467: data = 8'hca;
      17'd3468: data = 8'hf9;
      17'd3469: data = 8'h1b;
      17'd3470: data = 8'h05;
      17'd3471: data = 8'hf2;
      17'd3472: data = 8'hd6;
      17'd3473: data = 8'h16;
      17'd3474: data = 8'hfa;
      17'd3475: data = 8'hf9;
      17'd3476: data = 8'h0a;
      17'd3477: data = 8'hef;
      17'd3478: data = 8'h00;
      17'd3479: data = 8'he5;
      17'd3480: data = 8'h0d;
      17'd3481: data = 8'h1f;
      17'd3482: data = 8'hdc;
      17'd3483: data = 8'hde;
      17'd3484: data = 8'h15;
      17'd3485: data = 8'h15;
      17'd3486: data = 8'hf1;
      17'd3487: data = 8'hfc;
      17'd3488: data = 8'hf2;
      17'd3489: data = 8'h01;
      17'd3490: data = 8'h16;
      17'd3491: data = 8'h01;
      17'd3492: data = 8'he5;
      17'd3493: data = 8'h01;
      17'd3494: data = 8'h06;
      17'd3495: data = 8'h09;
      17'd3496: data = 8'h0d;
      17'd3497: data = 8'hce;
      17'd3498: data = 8'h05;
      17'd3499: data = 8'h23;
      17'd3500: data = 8'hdc;
      17'd3501: data = 8'hf9;
      17'd3502: data = 8'h26;
      17'd3503: data = 8'he7;
      17'd3504: data = 8'he2;
      17'd3505: data = 8'h13;
      17'd3506: data = 8'h11;
      17'd3507: data = 8'hf5;
      17'd3508: data = 8'hed;
      17'd3509: data = 8'h09;
      17'd3510: data = 8'hf5;
      17'd3511: data = 8'hfe;
      17'd3512: data = 8'h13;
      17'd3513: data = 8'he5;
      17'd3514: data = 8'hde;
      17'd3515: data = 8'h11;
      17'd3516: data = 8'h15;
      17'd3517: data = 8'hde;
      17'd3518: data = 8'hef;
      17'd3519: data = 8'h12;
      17'd3520: data = 8'h00;
      17'd3521: data = 8'hf2;
      17'd3522: data = 8'h01;
      17'd3523: data = 8'h05;
      17'd3524: data = 8'h06;
      17'd3525: data = 8'hf2;
      17'd3526: data = 8'hed;
      17'd3527: data = 8'h1a;
      17'd3528: data = 8'h0d;
      17'd3529: data = 8'hec;
      17'd3530: data = 8'hf9;
      17'd3531: data = 8'h09;
      17'd3532: data = 8'h1b;
      17'd3533: data = 8'h09;
      17'd3534: data = 8'hed;
      17'd3535: data = 8'h04;
      17'd3536: data = 8'h1a;
      17'd3537: data = 8'h1b;
      17'd3538: data = 8'he3;
      17'd3539: data = 8'h00;
      17'd3540: data = 8'h1a;
      17'd3541: data = 8'hfa;
      17'd3542: data = 8'hfe;
      17'd3543: data = 8'h11;
      17'd3544: data = 8'h05;
      17'd3545: data = 8'hec;
      17'd3546: data = 8'hfc;
      17'd3547: data = 8'h26;
      17'd3548: data = 8'h15;
      17'd3549: data = 8'heb;
      17'd3550: data = 8'h01;
      17'd3551: data = 8'h11;
      17'd3552: data = 8'h12;
      17'd3553: data = 8'h00;
      17'd3554: data = 8'hfc;
      17'd3555: data = 8'h0e;
      17'd3556: data = 8'h02;
      17'd3557: data = 8'hfa;
      17'd3558: data = 8'h04;
      17'd3559: data = 8'h15;
      17'd3560: data = 8'h00;
      17'd3561: data = 8'hfd;
      17'd3562: data = 8'h19;
      17'd3563: data = 8'hfc;
      17'd3564: data = 8'hf4;
      17'd3565: data = 8'h23;
      17'd3566: data = 8'h0a;
      17'd3567: data = 8'he7;
      17'd3568: data = 8'h05;
      17'd3569: data = 8'h09;
      17'd3570: data = 8'hfc;
      17'd3571: data = 8'hf9;
      17'd3572: data = 8'h02;
      17'd3573: data = 8'h0a;
      17'd3574: data = 8'hed;
      17'd3575: data = 8'hfd;
      17'd3576: data = 8'h15;
      17'd3577: data = 8'hf1;
      17'd3578: data = 8'h05;
      17'd3579: data = 8'h05;
      17'd3580: data = 8'heb;
      17'd3581: data = 8'hfa;
      17'd3582: data = 8'h15;
      17'd3583: data = 8'h04;
      17'd3584: data = 8'he0;
      17'd3585: data = 8'hfa;
      17'd3586: data = 8'h0e;
      17'd3587: data = 8'hfe;
      17'd3588: data = 8'hf9;
      17'd3589: data = 8'hfa;
      17'd3590: data = 8'hfc;
      17'd3591: data = 8'h00;
      17'd3592: data = 8'h06;
      17'd3593: data = 8'hfc;
      17'd3594: data = 8'hec;
      17'd3595: data = 8'h09;
      17'd3596: data = 8'h0e;
      17'd3597: data = 8'hf6;
      17'd3598: data = 8'hed;
      17'd3599: data = 8'h19;
      17'd3600: data = 8'h02;
      17'd3601: data = 8'hef;
      17'd3602: data = 8'h01;
      17'd3603: data = 8'h01;
      17'd3604: data = 8'h09;
      17'd3605: data = 8'he9;
      17'd3606: data = 8'h0e;
      17'd3607: data = 8'h06;
      17'd3608: data = 8'hd8;
      17'd3609: data = 8'h1b;
      17'd3610: data = 8'h16;
      17'd3611: data = 8'he3;
      17'd3612: data = 8'h05;
      17'd3613: data = 8'hf6;
      17'd3614: data = 8'h04;
      17'd3615: data = 8'h11;
      17'd3616: data = 8'heb;
      17'd3617: data = 8'hf2;
      17'd3618: data = 8'h01;
      17'd3619: data = 8'h0c;
      17'd3620: data = 8'hf1;
      17'd3621: data = 8'hfe;
      17'd3622: data = 8'h0e;
      17'd3623: data = 8'hec;
      17'd3624: data = 8'hef;
      17'd3625: data = 8'h09;
      17'd3626: data = 8'h09;
      17'd3627: data = 8'hef;
      17'd3628: data = 8'h04;
      17'd3629: data = 8'hef;
      17'd3630: data = 8'hf6;
      17'd3631: data = 8'h1c;
      17'd3632: data = 8'heb;
      17'd3633: data = 8'hfd;
      17'd3634: data = 8'h02;
      17'd3635: data = 8'hfc;
      17'd3636: data = 8'h1e;
      17'd3637: data = 8'hef;
      17'd3638: data = 8'he5;
      17'd3639: data = 8'h1a;
      17'd3640: data = 8'h19;
      17'd3641: data = 8'hec;
      17'd3642: data = 8'hd2;
      17'd3643: data = 8'h22;
      17'd3644: data = 8'h16;
      17'd3645: data = 8'hd8;
      17'd3646: data = 8'h0d;
      17'd3647: data = 8'h0d;
      17'd3648: data = 8'heb;
      17'd3649: data = 8'h1e;
      17'd3650: data = 8'h0a;
      17'd3651: data = 8'he3;
      17'd3652: data = 8'h16;
      17'd3653: data = 8'h09;
      17'd3654: data = 8'hef;
      17'd3655: data = 8'hf1;
      17'd3656: data = 8'h24;
      17'd3657: data = 8'h12;
      17'd3658: data = 8'hbb;
      17'd3659: data = 8'h01;
      17'd3660: data = 8'h31;
      17'd3661: data = 8'hf6;
      17'd3662: data = 8'he9;
      17'd3663: data = 8'h02;
      17'd3664: data = 8'hfa;
      17'd3665: data = 8'h0d;
      17'd3666: data = 8'h16;
      17'd3667: data = 8'he9;
      17'd3668: data = 8'hd2;
      17'd3669: data = 8'h15;
      17'd3670: data = 8'h31;
      17'd3671: data = 8'hd8;
      17'd3672: data = 8'hdb;
      17'd3673: data = 8'h12;
      17'd3674: data = 8'h12;
      17'd3675: data = 8'he7;
      17'd3676: data = 8'hed;
      17'd3677: data = 8'h0e;
      17'd3678: data = 8'hf9;
      17'd3679: data = 8'hf5;
      17'd3680: data = 8'hfa;
      17'd3681: data = 8'hfa;
      17'd3682: data = 8'h02;
      17'd3683: data = 8'h06;
      17'd3684: data = 8'hf2;
      17'd3685: data = 8'he2;
      17'd3686: data = 8'h06;
      17'd3687: data = 8'h22;
      17'd3688: data = 8'he2;
      17'd3689: data = 8'hd6;
      17'd3690: data = 8'h13;
      17'd3691: data = 8'h0c;
      17'd3692: data = 8'hd3;
      17'd3693: data = 8'hfc;
      17'd3694: data = 8'h24;
      17'd3695: data = 8'hda;
      17'd3696: data = 8'he9;
      17'd3697: data = 8'hfe;
      17'd3698: data = 8'h11;
      17'd3699: data = 8'h05;
      17'd3700: data = 8'hdb;
      17'd3701: data = 8'h04;
      17'd3702: data = 8'h0e;
      17'd3703: data = 8'hfe;
      17'd3704: data = 8'hed;
      17'd3705: data = 8'h02;
      17'd3706: data = 8'hf1;
      17'd3707: data = 8'h06;
      17'd3708: data = 8'h13;
      17'd3709: data = 8'hca;
      17'd3710: data = 8'h12;
      17'd3711: data = 8'h0d;
      17'd3712: data = 8'hdc;
      17'd3713: data = 8'h15;
      17'd3714: data = 8'h01;
      17'd3715: data = 8'hf5;
      17'd3716: data = 8'hf9;
      17'd3717: data = 8'hf5;
      17'd3718: data = 8'h1f;
      17'd3719: data = 8'hf5;
      17'd3720: data = 8'hf1;
      17'd3721: data = 8'h09;
      17'd3722: data = 8'hdb;
      17'd3723: data = 8'h0c;
      17'd3724: data = 8'h29;
      17'd3725: data = 8'hd5;
      17'd3726: data = 8'hd6;
      17'd3727: data = 8'h1f;
      17'd3728: data = 8'h0c;
      17'd3729: data = 8'he9;
      17'd3730: data = 8'hf5;
      17'd3731: data = 8'h0c;
      17'd3732: data = 8'h0d;
      17'd3733: data = 8'he4;
      17'd3734: data = 8'hed;
      17'd3735: data = 8'h16;
      17'd3736: data = 8'hfe;
      17'd3737: data = 8'hfd;
      17'd3738: data = 8'hf4;
      17'd3739: data = 8'he5;
      17'd3740: data = 8'h1c;
      17'd3741: data = 8'h13;
      17'd3742: data = 8'he0;
      17'd3743: data = 8'hfe;
      17'd3744: data = 8'h23;
      17'd3745: data = 8'hf5;
      17'd3746: data = 8'hf4;
      17'd3747: data = 8'h1b;
      17'd3748: data = 8'h01;
      17'd3749: data = 8'hfc;
      17'd3750: data = 8'hfc;
      17'd3751: data = 8'h04;
      17'd3752: data = 8'h12;
      17'd3753: data = 8'he7;
      17'd3754: data = 8'h00;
      17'd3755: data = 8'h0d;
      17'd3756: data = 8'hf6;
      17'd3757: data = 8'h1e;
      17'd3758: data = 8'hf9;
      17'd3759: data = 8'hde;
      17'd3760: data = 8'h1b;
      17'd3761: data = 8'h1a;
      17'd3762: data = 8'he5;
      17'd3763: data = 8'hec;
      17'd3764: data = 8'h15;
      17'd3765: data = 8'h13;
      17'd3766: data = 8'hec;
      17'd3767: data = 8'hfa;
      17'd3768: data = 8'h16;
      17'd3769: data = 8'hf4;
      17'd3770: data = 8'h04;
      17'd3771: data = 8'h1a;
      17'd3772: data = 8'hfe;
      17'd3773: data = 8'hfc;
      17'd3774: data = 8'h05;
      17'd3775: data = 8'h0a;
      17'd3776: data = 8'h0c;
      17'd3777: data = 8'h04;
      17'd3778: data = 8'h00;
      17'd3779: data = 8'hfc;
      17'd3780: data = 8'h05;
      17'd3781: data = 8'h0d;
      17'd3782: data = 8'h04;
      17'd3783: data = 8'hf5;
      17'd3784: data = 8'h09;
      17'd3785: data = 8'h26;
      17'd3786: data = 8'he0;
      17'd3787: data = 8'heb;
      17'd3788: data = 8'h31;
      17'd3789: data = 8'h00;
      17'd3790: data = 8'hf2;
      17'd3791: data = 8'h09;
      17'd3792: data = 8'hf4;
      17'd3793: data = 8'hfc;
      17'd3794: data = 8'h19;
      17'd3795: data = 8'h04;
      17'd3796: data = 8'hed;
      17'd3797: data = 8'hf9;
      17'd3798: data = 8'h02;
      17'd3799: data = 8'h0c;
      17'd3800: data = 8'h0a;
      17'd3801: data = 8'hf5;
      17'd3802: data = 8'hed;
      17'd3803: data = 8'h0e;
      17'd3804: data = 8'h1e;
      17'd3805: data = 8'h00;
      17'd3806: data = 8'he0;
      17'd3807: data = 8'h06;
      17'd3808: data = 8'h19;
      17'd3809: data = 8'h06;
      17'd3810: data = 8'heb;
      17'd3811: data = 8'hec;
      17'd3812: data = 8'h26;
      17'd3813: data = 8'h02;
      17'd3814: data = 8'hf1;
      17'd3815: data = 8'h00;
      17'd3816: data = 8'h0a;
      17'd3817: data = 8'hfe;
      17'd3818: data = 8'hf4;
      17'd3819: data = 8'h15;
      17'd3820: data = 8'h04;
      17'd3821: data = 8'heb;
      17'd3822: data = 8'hf4;
      17'd3823: data = 8'h0e;
      17'd3824: data = 8'h0e;
      17'd3825: data = 8'hf4;
      17'd3826: data = 8'hfa;
      17'd3827: data = 8'hf6;
      17'd3828: data = 8'h00;
      17'd3829: data = 8'h27;
      17'd3830: data = 8'hf2;
      17'd3831: data = 8'hd5;
      17'd3832: data = 8'h1e;
      17'd3833: data = 8'h13;
      17'd3834: data = 8'he4;
      17'd3835: data = 8'hf1;
      17'd3836: data = 8'h0d;
      17'd3837: data = 8'hf5;
      17'd3838: data = 8'hfd;
      17'd3839: data = 8'h1b;
      17'd3840: data = 8'he7;
      17'd3841: data = 8'hd3;
      17'd3842: data = 8'h40;
      17'd3843: data = 8'h0c;
      17'd3844: data = 8'hbd;
      17'd3845: data = 8'h1e;
      17'd3846: data = 8'h1b;
      17'd3847: data = 8'he0;
      17'd3848: data = 8'hfa;
      17'd3849: data = 8'h1c;
      17'd3850: data = 8'h04;
      17'd3851: data = 8'hc9;
      17'd3852: data = 8'h05;
      17'd3853: data = 8'h40;
      17'd3854: data = 8'he5;
      17'd3855: data = 8'he0;
      17'd3856: data = 8'h1c;
      17'd3857: data = 8'h00;
      17'd3858: data = 8'hfe;
      17'd3859: data = 8'h2d;
      17'd3860: data = 8'hda;
      17'd3861: data = 8'hd8;
      17'd3862: data = 8'h40;
      17'd3863: data = 8'h0a;
      17'd3864: data = 8'hbc;
      17'd3865: data = 8'h05;
      17'd3866: data = 8'h42;
      17'd3867: data = 8'hdc;
      17'd3868: data = 8'hd1;
      17'd3869: data = 8'h31;
      17'd3870: data = 8'h19;
      17'd3871: data = 8'hd3;
      17'd3872: data = 8'h06;
      17'd3873: data = 8'h01;
      17'd3874: data = 8'hf9;
      17'd3875: data = 8'h1c;
      17'd3876: data = 8'he0;
      17'd3877: data = 8'he9;
      17'd3878: data = 8'h0e;
      17'd3879: data = 8'h12;
      17'd3880: data = 8'hef;
      17'd3881: data = 8'hd2;
      17'd3882: data = 8'h1a;
      17'd3883: data = 8'h1a;
      17'd3884: data = 8'hdb;
      17'd3885: data = 8'hf5;
      17'd3886: data = 8'h05;
      17'd3887: data = 8'h04;
      17'd3888: data = 8'hfe;
      17'd3889: data = 8'hdc;
      17'd3890: data = 8'h01;
      17'd3891: data = 8'h19;
      17'd3892: data = 8'hf2;
      17'd3893: data = 8'hdb;
      17'd3894: data = 8'hf4;
      17'd3895: data = 8'h16;
      17'd3896: data = 8'h16;
      17'd3897: data = 8'hd3;
      17'd3898: data = 8'hf1;
      17'd3899: data = 8'h19;
      17'd3900: data = 8'hf2;
      17'd3901: data = 8'hfc;
      17'd3902: data = 8'hf5;
      17'd3903: data = 8'h06;
      17'd3904: data = 8'hf9;
      17'd3905: data = 8'he9;
      17'd3906: data = 8'hf6;
      17'd3907: data = 8'h01;
      17'd3908: data = 8'h22;
      17'd3909: data = 8'hf2;
      17'd3910: data = 8'hc9;
      17'd3911: data = 8'h0c;
      17'd3912: data = 8'h29;
      17'd3913: data = 8'hef;
      17'd3914: data = 8'hd8;
      17'd3915: data = 8'hfd;
      17'd3916: data = 8'h1b;
      17'd3917: data = 8'hf2;
      17'd3918: data = 8'he3;
      17'd3919: data = 8'h0c;
      17'd3920: data = 8'hef;
      17'd3921: data = 8'hf4;
      17'd3922: data = 8'h22;
      17'd3923: data = 8'he9;
      17'd3924: data = 8'he5;
      17'd3925: data = 8'h1a;
      17'd3926: data = 8'he4;
      17'd3927: data = 8'he4;
      17'd3928: data = 8'h35;
      17'd3929: data = 8'hef;
      17'd3930: data = 8'hc5;
      17'd3931: data = 8'h1e;
      17'd3932: data = 8'h0e;
      17'd3933: data = 8'hed;
      17'd3934: data = 8'hf9;
      17'd3935: data = 8'hfd;
      17'd3936: data = 8'hf9;
      17'd3937: data = 8'hf1;
      17'd3938: data = 8'h11;
      17'd3939: data = 8'h00;
      17'd3940: data = 8'heb;
      17'd3941: data = 8'hfc;
      17'd3942: data = 8'hf2;
      17'd3943: data = 8'h09;
      17'd3944: data = 8'h1a;
      17'd3945: data = 8'hef;
      17'd3946: data = 8'hd2;
      17'd3947: data = 8'h12;
      17'd3948: data = 8'h27;
      17'd3949: data = 8'hfa;
      17'd3950: data = 8'hc6;
      17'd3951: data = 8'h1c;
      17'd3952: data = 8'h19;
      17'd3953: data = 8'hc5;
      17'd3954: data = 8'h1b;
      17'd3955: data = 8'h04;
      17'd3956: data = 8'hf5;
      17'd3957: data = 8'h09;
      17'd3958: data = 8'hf9;
      17'd3959: data = 8'hfe;
      17'd3960: data = 8'h00;
      17'd3961: data = 8'h15;
      17'd3962: data = 8'h02;
      17'd3963: data = 8'hda;
      17'd3964: data = 8'h04;
      17'd3965: data = 8'h1e;
      17'd3966: data = 8'hf1;
      17'd3967: data = 8'hf2;
      17'd3968: data = 8'hfd;
      17'd3969: data = 8'h0a;
      17'd3970: data = 8'hfd;
      17'd3971: data = 8'he4;
      17'd3972: data = 8'h04;
      17'd3973: data = 8'h0a;
      17'd3974: data = 8'h01;
      17'd3975: data = 8'hf2;
      17'd3976: data = 8'he2;
      17'd3977: data = 8'h24;
      17'd3978: data = 8'h05;
      17'd3979: data = 8'hcb;
      17'd3980: data = 8'h1a;
      17'd3981: data = 8'h09;
      17'd3982: data = 8'hda;
      17'd3983: data = 8'h06;
      17'd3984: data = 8'h11;
      17'd3985: data = 8'hfa;
      17'd3986: data = 8'hef;
      17'd3987: data = 8'hf6;
      17'd3988: data = 8'h13;
      17'd3989: data = 8'h09;
      17'd3990: data = 8'hf1;
      17'd3991: data = 8'he7;
      17'd3992: data = 8'h0c;
      17'd3993: data = 8'h1e;
      17'd3994: data = 8'hf4;
      17'd3995: data = 8'heb;
      17'd3996: data = 8'hf9;
      17'd3997: data = 8'h29;
      17'd3998: data = 8'h04;
      17'd3999: data = 8'hd3;
      17'd4000: data = 8'h0d;
      17'd4001: data = 8'h1f;
      17'd4002: data = 8'hfd;
      17'd4003: data = 8'hde;
      17'd4004: data = 8'hf9;
      17'd4005: data = 8'h26;
      17'd4006: data = 8'h13;
      17'd4007: data = 8'hda;
      17'd4008: data = 8'hfc;
      17'd4009: data = 8'h0e;
      17'd4010: data = 8'h16;
      17'd4011: data = 8'h0c;
      17'd4012: data = 8'hda;
      17'd4013: data = 8'h04;
      17'd4014: data = 8'h1e;
      17'd4015: data = 8'hf5;
      17'd4016: data = 8'hfd;
      17'd4017: data = 8'hfd;
      17'd4018: data = 8'h00;
      17'd4019: data = 8'h0e;
      17'd4020: data = 8'hec;
      17'd4021: data = 8'h06;
      17'd4022: data = 8'h15;
      17'd4023: data = 8'hf5;
      17'd4024: data = 8'h00;
      17'd4025: data = 8'hfd;
      17'd4026: data = 8'h12;
      17'd4027: data = 8'h11;
      17'd4028: data = 8'hde;
      17'd4029: data = 8'hfc;
      17'd4030: data = 8'h1b;
      17'd4031: data = 8'h0c;
      17'd4032: data = 8'hde;
      17'd4033: data = 8'hf6;
      17'd4034: data = 8'h27;
      17'd4035: data = 8'hef;
      17'd4036: data = 8'hfd;
      17'd4037: data = 8'h0a;
      17'd4038: data = 8'h00;
      17'd4039: data = 8'hfa;
      17'd4040: data = 8'hf5;
      17'd4041: data = 8'h16;
      17'd4042: data = 8'h01;
      17'd4043: data = 8'he4;
      17'd4044: data = 8'h09;
      17'd4045: data = 8'h09;
      17'd4046: data = 8'hf6;
      17'd4047: data = 8'h12;
      17'd4048: data = 8'hf6;
      17'd4049: data = 8'he4;
      17'd4050: data = 8'h1e;
      17'd4051: data = 8'h1e;
      17'd4052: data = 8'hd6;
      17'd4053: data = 8'he5;
      17'd4054: data = 8'h2b;
      17'd4055: data = 8'h1a;
      17'd4056: data = 8'hda;
      17'd4057: data = 8'hdb;
      17'd4058: data = 8'h1c;
      17'd4059: data = 8'h36;
      17'd4060: data = 8'hdb;
      17'd4061: data = 8'hdc;
      17'd4062: data = 8'h23;
      17'd4063: data = 8'h1f;
      17'd4064: data = 8'h09;
      17'd4065: data = 8'he4;
      17'd4066: data = 8'h00;
      17'd4067: data = 8'h31;
      17'd4068: data = 8'h01;
      17'd4069: data = 8'he0;
      17'd4070: data = 8'h13;
      17'd4071: data = 8'hfd;
      17'd4072: data = 8'h04;
      17'd4073: data = 8'h1a;
      17'd4074: data = 8'h01;
      17'd4075: data = 8'hef;
      17'd4076: data = 8'hf4;
      17'd4077: data = 8'h1c;
      17'd4078: data = 8'h16;
      17'd4079: data = 8'he9;
      17'd4080: data = 8'h06;
      17'd4081: data = 8'h05;
      17'd4082: data = 8'hef;
      17'd4083: data = 8'h27;
      17'd4084: data = 8'hf6;
      17'd4085: data = 8'hf2;
      17'd4086: data = 8'h04;
      17'd4087: data = 8'hfc;
      17'd4088: data = 8'h0e;
      17'd4089: data = 8'hfe;
      17'd4090: data = 8'h00;
      17'd4091: data = 8'he9;
      17'd4092: data = 8'h04;
      17'd4093: data = 8'h19;
      17'd4094: data = 8'he3;
      17'd4095: data = 8'hf6;
      17'd4096: data = 8'h0d;
      17'd4097: data = 8'hf6;
      17'd4098: data = 8'hf2;
      17'd4099: data = 8'hfe;
      17'd4100: data = 8'h15;
      17'd4101: data = 8'hdc;
      17'd4102: data = 8'heb;
      17'd4103: data = 8'h31;
      17'd4104: data = 8'hfa;
      17'd4105: data = 8'hed;
      17'd4106: data = 8'hf2;
      17'd4107: data = 8'hfd;
      17'd4108: data = 8'h1a;
      17'd4109: data = 8'h01;
      17'd4110: data = 8'he3;
      17'd4111: data = 8'h05;
      17'd4112: data = 8'h1a;
      17'd4113: data = 8'hfa;
      17'd4114: data = 8'hf9;
      17'd4115: data = 8'h00;
      17'd4116: data = 8'h1f;
      17'd4117: data = 8'hfe;
      17'd4118: data = 8'hdb;
      17'd4119: data = 8'h0d;
      17'd4120: data = 8'h1c;
      17'd4121: data = 8'hfe;
      17'd4122: data = 8'hfd;
      17'd4123: data = 8'hf5;
      17'd4124: data = 8'hf6;
      17'd4125: data = 8'h39;
      17'd4126: data = 8'hf1;
      17'd4127: data = 8'hda;
      17'd4128: data = 8'h27;
      17'd4129: data = 8'h04;
      17'd4130: data = 8'hed;
      17'd4131: data = 8'hf6;
      17'd4132: data = 8'h13;
      17'd4133: data = 8'h0e;
      17'd4134: data = 8'hde;
      17'd4135: data = 8'hf6;
      17'd4136: data = 8'h1e;
      17'd4137: data = 8'hf9;
      17'd4138: data = 8'h0a;
      17'd4139: data = 8'hf5;
      17'd4140: data = 8'hde;
      17'd4141: data = 8'h24;
      17'd4142: data = 8'hf2;
      17'd4143: data = 8'h04;
      17'd4144: data = 8'hf9;
      17'd4145: data = 8'hd6;
      17'd4146: data = 8'h27;
      17'd4147: data = 8'hec;
      17'd4148: data = 8'hf1;
      17'd4149: data = 8'h0c;
      17'd4150: data = 8'he9;
      17'd4151: data = 8'h09;
      17'd4152: data = 8'h05;
      17'd4153: data = 8'hdb;
      17'd4154: data = 8'h09;
      17'd4155: data = 8'h19;
      17'd4156: data = 8'he3;
      17'd4157: data = 8'hed;
      17'd4158: data = 8'h0e;
      17'd4159: data = 8'h00;
      17'd4160: data = 8'heb;
      17'd4161: data = 8'hef;
      17'd4162: data = 8'h0a;
      17'd4163: data = 8'h24;
      17'd4164: data = 8'hdb;
      17'd4165: data = 8'h05;
      17'd4166: data = 8'h04;
      17'd4167: data = 8'h01;
      17'd4168: data = 8'h1e;
      17'd4169: data = 8'he9;
      17'd4170: data = 8'hf5;
      17'd4171: data = 8'h13;
      17'd4172: data = 8'h0a;
      17'd4173: data = 8'hf9;
      17'd4174: data = 8'h05;
      17'd4175: data = 8'h01;
      17'd4176: data = 8'h0c;
      17'd4177: data = 8'h05;
      17'd4178: data = 8'hfe;
      17'd4179: data = 8'h1b;
      17'd4180: data = 8'hf9;
      17'd4181: data = 8'he9;
      17'd4182: data = 8'h13;
      17'd4183: data = 8'h06;
      17'd4184: data = 8'hfe;
      17'd4185: data = 8'heb;
      17'd4186: data = 8'hf4;
      17'd4187: data = 8'h2d;
      17'd4188: data = 8'hf5;
      17'd4189: data = 8'hf1;
      17'd4190: data = 8'hfd;
      17'd4191: data = 8'hfc;
      17'd4192: data = 8'h22;
      17'd4193: data = 8'hfe;
      17'd4194: data = 8'he3;
      17'd4195: data = 8'hf6;
      17'd4196: data = 8'h1a;
      17'd4197: data = 8'hfa;
      17'd4198: data = 8'hde;
      17'd4199: data = 8'h01;
      17'd4200: data = 8'h09;
      17'd4201: data = 8'h01;
      17'd4202: data = 8'hef;
      17'd4203: data = 8'h02;
      17'd4204: data = 8'hfd;
      17'd4205: data = 8'hfd;
      17'd4206: data = 8'h15;
      17'd4207: data = 8'hde;
      17'd4208: data = 8'hf9;
      17'd4209: data = 8'h16;
      17'd4210: data = 8'h00;
      17'd4211: data = 8'he7;
      17'd4212: data = 8'he9;
      17'd4213: data = 8'h1a;
      17'd4214: data = 8'h0e;
      17'd4215: data = 8'he2;
      17'd4216: data = 8'he9;
      17'd4217: data = 8'h29;
      17'd4218: data = 8'h09;
      17'd4219: data = 8'hde;
      17'd4220: data = 8'h00;
      17'd4221: data = 8'h0c;
      17'd4222: data = 8'hfc;
      17'd4223: data = 8'hfc;
      17'd4224: data = 8'h04;
      17'd4225: data = 8'hfc;
      17'd4226: data = 8'hf1;
      17'd4227: data = 8'h01;
      17'd4228: data = 8'h13;
      17'd4229: data = 8'hfa;
      17'd4230: data = 8'hfe;
      17'd4231: data = 8'h01;
      17'd4232: data = 8'h15;
      17'd4233: data = 8'hed;
      17'd4234: data = 8'heb;
      17'd4235: data = 8'h31;
      17'd4236: data = 8'hfc;
      17'd4237: data = 8'hdc;
      17'd4238: data = 8'hfe;
      17'd4239: data = 8'h31;
      17'd4240: data = 8'he9;
      17'd4241: data = 8'hef;
      17'd4242: data = 8'h16;
      17'd4243: data = 8'h05;
      17'd4244: data = 8'h0d;
      17'd4245: data = 8'hdb;
      17'd4246: data = 8'h0d;
      17'd4247: data = 8'h0c;
      17'd4248: data = 8'h00;
      17'd4249: data = 8'hfa;
      17'd4250: data = 8'he2;
      17'd4251: data = 8'h16;
      17'd4252: data = 8'h0e;
      17'd4253: data = 8'he2;
      17'd4254: data = 8'hfd;
      17'd4255: data = 8'h01;
      17'd4256: data = 8'h15;
      17'd4257: data = 8'hf5;
      17'd4258: data = 8'hd6;
      17'd4259: data = 8'h3a;
      17'd4260: data = 8'hfe;
      17'd4261: data = 8'hc1;
      17'd4262: data = 8'h12;
      17'd4263: data = 8'h1b;
      17'd4264: data = 8'h0a;
      17'd4265: data = 8'hd6;
      17'd4266: data = 8'he3;
      17'd4267: data = 8'h2d;
      17'd4268: data = 8'h02;
      17'd4269: data = 8'hfa;
      17'd4270: data = 8'hf9;
      17'd4271: data = 8'hf6;
      17'd4272: data = 8'h12;
      17'd4273: data = 8'h0d;
      17'd4274: data = 8'hf9;
      17'd4275: data = 8'hef;
      17'd4276: data = 8'h1e;
      17'd4277: data = 8'hf9;
      17'd4278: data = 8'hec;
      17'd4279: data = 8'h1a;
      17'd4280: data = 8'h0e;
      17'd4281: data = 8'hec;
      17'd4282: data = 8'hf6;
      17'd4283: data = 8'h24;
      17'd4284: data = 8'hfa;
      17'd4285: data = 8'he4;
      17'd4286: data = 8'h24;
      17'd4287: data = 8'h04;
      17'd4288: data = 8'he5;
      17'd4289: data = 8'h19;
      17'd4290: data = 8'h09;
      17'd4291: data = 8'hf2;
      17'd4292: data = 8'h05;
      17'd4293: data = 8'h0a;
      17'd4294: data = 8'hfd;
      17'd4295: data = 8'h02;
      17'd4296: data = 8'h06;
      17'd4297: data = 8'hf5;
      17'd4298: data = 8'h01;
      17'd4299: data = 8'h13;
      17'd4300: data = 8'heb;
      17'd4301: data = 8'h0a;
      17'd4302: data = 8'h15;
      17'd4303: data = 8'hf6;
      17'd4304: data = 8'hed;
      17'd4305: data = 8'h0a;
      17'd4306: data = 8'h1e;
      17'd4307: data = 8'he0;
      17'd4308: data = 8'heb;
      17'd4309: data = 8'h23;
      17'd4310: data = 8'hfc;
      17'd4311: data = 8'hd2;
      17'd4312: data = 8'h1a;
      17'd4313: data = 8'h15;
      17'd4314: data = 8'hd1;
      17'd4315: data = 8'hfd;
      17'd4316: data = 8'h2c;
      17'd4317: data = 8'hec;
      17'd4318: data = 8'hde;
      17'd4319: data = 8'h2b;
      17'd4320: data = 8'hfa;
      17'd4321: data = 8'he0;
      17'd4322: data = 8'h23;
      17'd4323: data = 8'hfd;
      17'd4324: data = 8'hde;
      17'd4325: data = 8'h0e;
      17'd4326: data = 8'h06;
      17'd4327: data = 8'hf9;
      17'd4328: data = 8'hfa;
      17'd4329: data = 8'hf4;
      17'd4330: data = 8'h19;
      17'd4331: data = 8'hfa;
      17'd4332: data = 8'hf4;
      17'd4333: data = 8'h26;
      17'd4334: data = 8'hfd;
      17'd4335: data = 8'he5;
      17'd4336: data = 8'h1b;
      17'd4337: data = 8'hfc;
      17'd4338: data = 8'hfc;
      17'd4339: data = 8'h0d;
      17'd4340: data = 8'hfd;
      17'd4341: data = 8'h0c;
      17'd4342: data = 8'he9;
      17'd4343: data = 8'h13;
      17'd4344: data = 8'h0a;
      17'd4345: data = 8'he7;
      17'd4346: data = 8'h19;
      17'd4347: data = 8'h02;
      17'd4348: data = 8'he4;
      17'd4349: data = 8'h12;
      17'd4350: data = 8'hf9;
      17'd4351: data = 8'h00;
      17'd4352: data = 8'h0c;
      17'd4353: data = 8'he0;
      17'd4354: data = 8'h0c;
      17'd4355: data = 8'hf9;
      17'd4356: data = 8'h0d;
      17'd4357: data = 8'h05;
      17'd4358: data = 8'he2;
      17'd4359: data = 8'hfc;
      17'd4360: data = 8'h16;
      17'd4361: data = 8'hec;
      17'd4362: data = 8'h0a;
      17'd4363: data = 8'h0d;
      17'd4364: data = 8'hce;
      17'd4365: data = 8'h00;
      17'd4366: data = 8'h1c;
      17'd4367: data = 8'h0e;
      17'd4368: data = 8'hc5;
      17'd4369: data = 8'hfe;
      17'd4370: data = 8'h16;
      17'd4371: data = 8'hf2;
      17'd4372: data = 8'h04;
      17'd4373: data = 8'h02;
      17'd4374: data = 8'he3;
      17'd4375: data = 8'hfa;
      17'd4376: data = 8'h1f;
      17'd4377: data = 8'hf2;
      17'd4378: data = 8'h06;
      17'd4379: data = 8'hed;
      17'd4380: data = 8'he5;
      17'd4381: data = 8'h2c;
      17'd4382: data = 8'h05;
      17'd4383: data = 8'he4;
      17'd4384: data = 8'h05;
      17'd4385: data = 8'hf4;
      17'd4386: data = 8'h0c;
      17'd4387: data = 8'h22;
      17'd4388: data = 8'hd5;
      17'd4389: data = 8'hec;
      17'd4390: data = 8'h2b;
      17'd4391: data = 8'h0a;
      17'd4392: data = 8'he9;
      17'd4393: data = 8'hf9;
      17'd4394: data = 8'h05;
      17'd4395: data = 8'h16;
      17'd4396: data = 8'hf4;
      17'd4397: data = 8'hfc;
      17'd4398: data = 8'h02;
      17'd4399: data = 8'he7;
      17'd4400: data = 8'h11;
      17'd4401: data = 8'h0d;
      17'd4402: data = 8'hf5;
      17'd4403: data = 8'hed;
      17'd4404: data = 8'h00;
      17'd4405: data = 8'h00;
      17'd4406: data = 8'h04;
      17'd4407: data = 8'h13;
      17'd4408: data = 8'he9;
      17'd4409: data = 8'he0;
      17'd4410: data = 8'hfc;
      17'd4411: data = 8'h29;
      17'd4412: data = 8'h02;
      17'd4413: data = 8'hcd;
      17'd4414: data = 8'hfd;
      17'd4415: data = 8'h0a;
      17'd4416: data = 8'h0d;
      17'd4417: data = 8'h00;
      17'd4418: data = 8'hec;
      17'd4419: data = 8'hf1;
      17'd4420: data = 8'h0a;
      17'd4421: data = 8'h05;
      17'd4422: data = 8'hfe;
      17'd4423: data = 8'hfc;
      17'd4424: data = 8'hf5;
      17'd4425: data = 8'h01;
      17'd4426: data = 8'hf6;
      17'd4427: data = 8'h16;
      17'd4428: data = 8'h0a;
      17'd4429: data = 8'hda;
      17'd4430: data = 8'h02;
      17'd4431: data = 8'h2b;
      17'd4432: data = 8'h05;
      17'd4433: data = 8'hda;
      17'd4434: data = 8'h02;
      17'd4435: data = 8'h1b;
      17'd4436: data = 8'hfe;
      17'd4437: data = 8'h05;
      17'd4438: data = 8'heb;
      17'd4439: data = 8'hfa;
      17'd4440: data = 8'h0c;
      17'd4441: data = 8'h0a;
      17'd4442: data = 8'h0e;
      17'd4443: data = 8'hd6;
      17'd4444: data = 8'h00;
      17'd4445: data = 8'h1c;
      17'd4446: data = 8'hf2;
      17'd4447: data = 8'hfd;
      17'd4448: data = 8'h00;
      17'd4449: data = 8'h09;
      17'd4450: data = 8'h0e;
      17'd4451: data = 8'hd3;
      17'd4452: data = 8'h0c;
      17'd4453: data = 8'h1e;
      17'd4454: data = 8'he2;
      17'd4455: data = 8'hfe;
      17'd4456: data = 8'h04;
      17'd4457: data = 8'hfd;
      17'd4458: data = 8'h06;
      17'd4459: data = 8'hed;
      17'd4460: data = 8'h00;
      17'd4461: data = 8'h19;
      17'd4462: data = 8'he4;
      17'd4463: data = 8'hf5;
      17'd4464: data = 8'h09;
      17'd4465: data = 8'h0c;
      17'd4466: data = 8'hf2;
      17'd4467: data = 8'hf5;
      17'd4468: data = 8'hfc;
      17'd4469: data = 8'h02;
      17'd4470: data = 8'h05;
      17'd4471: data = 8'hed;
      17'd4472: data = 8'h06;
      17'd4473: data = 8'hf2;
      17'd4474: data = 8'hf5;
      17'd4475: data = 8'h1e;
      17'd4476: data = 8'hfe;
      17'd4477: data = 8'hd3;
      17'd4478: data = 8'h15;
      17'd4479: data = 8'h15;
      17'd4480: data = 8'he5;
      17'd4481: data = 8'hfc;
      17'd4482: data = 8'h06;
      17'd4483: data = 8'h01;
      17'd4484: data = 8'hfc;
      17'd4485: data = 8'h00;
      17'd4486: data = 8'h05;
      17'd4487: data = 8'h0c;
      17'd4488: data = 8'hf4;
      17'd4489: data = 8'hfd;
      17'd4490: data = 8'h15;
      17'd4491: data = 8'hf4;
      17'd4492: data = 8'hef;
      17'd4493: data = 8'h1a;
      17'd4494: data = 8'h0c;
      17'd4495: data = 8'he3;
      17'd4496: data = 8'hf2;
      17'd4497: data = 8'h15;
      17'd4498: data = 8'h15;
      17'd4499: data = 8'hf6;
      17'd4500: data = 8'hed;
      17'd4501: data = 8'h0c;
      17'd4502: data = 8'h0a;
      17'd4503: data = 8'hfa;
      17'd4504: data = 8'he7;
      17'd4505: data = 8'h19;
      17'd4506: data = 8'h04;
      17'd4507: data = 8'he7;
      17'd4508: data = 8'h12;
      17'd4509: data = 8'hec;
      17'd4510: data = 8'h06;
      17'd4511: data = 8'h0e;
      17'd4512: data = 8'h0c;
      17'd4513: data = 8'hfc;
      17'd4514: data = 8'he0;
      17'd4515: data = 8'h29;
      17'd4516: data = 8'h01;
      17'd4517: data = 8'hcd;
      17'd4518: data = 8'h23;
      17'd4519: data = 8'h0a;
      17'd4520: data = 8'hef;
      17'd4521: data = 8'hec;
      17'd4522: data = 8'hfe;
      17'd4523: data = 8'h1a;
      17'd4524: data = 8'hed;
      17'd4525: data = 8'h12;
      17'd4526: data = 8'hec;
      17'd4527: data = 8'hed;
      17'd4528: data = 8'h2b;
      17'd4529: data = 8'heb;
      17'd4530: data = 8'hf4;
      17'd4531: data = 8'h13;
      17'd4532: data = 8'hf6;
      17'd4533: data = 8'hfa;
      17'd4534: data = 8'hfa;
      17'd4535: data = 8'hfc;
      17'd4536: data = 8'h19;
      17'd4537: data = 8'h09;
      17'd4538: data = 8'hdb;
      17'd4539: data = 8'hfa;
      17'd4540: data = 8'h19;
      17'd4541: data = 8'h1c;
      17'd4542: data = 8'hf5;
      17'd4543: data = 8'hd2;
      17'd4544: data = 8'h1c;
      17'd4545: data = 8'h0a;
      17'd4546: data = 8'hfe;
      17'd4547: data = 8'h00;
      17'd4548: data = 8'hfa;
      17'd4549: data = 8'h0a;
      17'd4550: data = 8'hed;
      17'd4551: data = 8'h1b;
      17'd4552: data = 8'h0e;
      17'd4553: data = 8'hdb;
      17'd4554: data = 8'h12;
      17'd4555: data = 8'h12;
      17'd4556: data = 8'he9;
      17'd4557: data = 8'h09;
      17'd4558: data = 8'h05;
      17'd4559: data = 8'he5;
      17'd4560: data = 8'h1f;
      17'd4561: data = 8'h16;
      17'd4562: data = 8'hcd;
      17'd4563: data = 8'h00;
      17'd4564: data = 8'h1c;
      17'd4565: data = 8'h00;
      17'd4566: data = 8'hef;
      17'd4567: data = 8'hef;
      17'd4568: data = 8'h0d;
      17'd4569: data = 8'h09;
      17'd4570: data = 8'hed;
      17'd4571: data = 8'hef;
      17'd4572: data = 8'h0c;
      17'd4573: data = 8'h0a;
      17'd4574: data = 8'hed;
      17'd4575: data = 8'hef;
      17'd4576: data = 8'hf2;
      17'd4577: data = 8'h29;
      17'd4578: data = 8'h15;
      17'd4579: data = 8'hab;
      17'd4580: data = 8'h01;
      17'd4581: data = 8'h42;
      17'd4582: data = 8'hd1;
      17'd4583: data = 8'he9;
      17'd4584: data = 8'h23;
      17'd4585: data = 8'he7;
      17'd4586: data = 8'he9;
      17'd4587: data = 8'h02;
      17'd4588: data = 8'h1c;
      17'd4589: data = 8'hf6;
      17'd4590: data = 8'hde;
      17'd4591: data = 8'h0e;
      17'd4592: data = 8'h05;
      17'd4593: data = 8'hfc;
      17'd4594: data = 8'he2;
      17'd4595: data = 8'h13;
      17'd4596: data = 8'h1a;
      17'd4597: data = 8'hd2;
      17'd4598: data = 8'h1c;
      17'd4599: data = 8'hf9;
      17'd4600: data = 8'he4;
      17'd4601: data = 8'h2b;
      17'd4602: data = 8'hfe;
      17'd4603: data = 8'he7;
      17'd4604: data = 8'h02;
      17'd4605: data = 8'hf4;
      17'd4606: data = 8'h00;
      17'd4607: data = 8'h34;
      17'd4608: data = 8'he3;
      17'd4609: data = 8'he9;
      17'd4610: data = 8'h0d;
      17'd4611: data = 8'hfe;
      17'd4612: data = 8'h1f;
      17'd4613: data = 8'he7;
      17'd4614: data = 8'hec;
      17'd4615: data = 8'h15;
      17'd4616: data = 8'h04;
      17'd4617: data = 8'heb;
      17'd4618: data = 8'h1a;
      17'd4619: data = 8'hfe;
      17'd4620: data = 8'hc6;
      17'd4621: data = 8'h1c;
      17'd4622: data = 8'h15;
      17'd4623: data = 8'hfa;
      17'd4624: data = 8'he5;
      17'd4625: data = 8'heb;
      17'd4626: data = 8'h1f;
      17'd4627: data = 8'hfe;
      17'd4628: data = 8'h01;
      17'd4629: data = 8'hf1;
      17'd4630: data = 8'hde;
      17'd4631: data = 8'h1a;
      17'd4632: data = 8'h11;
      17'd4633: data = 8'he2;
      17'd4634: data = 8'hec;
      17'd4635: data = 8'h0e;
      17'd4636: data = 8'h04;
      17'd4637: data = 8'hec;
      17'd4638: data = 8'h06;
      17'd4639: data = 8'h13;
      17'd4640: data = 8'hed;
      17'd4641: data = 8'hf5;
      17'd4642: data = 8'h0e;
      17'd4643: data = 8'hf1;
      17'd4644: data = 8'hfc;
      17'd4645: data = 8'h35;
      17'd4646: data = 8'he2;
      17'd4647: data = 8'hcd;
      17'd4648: data = 8'h3a;
      17'd4649: data = 8'h0a;
      17'd4650: data = 8'hce;
      17'd4651: data = 8'h12;
      17'd4652: data = 8'h1f;
      17'd4653: data = 8'he7;
      17'd4654: data = 8'hef;
      17'd4655: data = 8'h11;
      17'd4656: data = 8'h1b;
      17'd4657: data = 8'hdb;
      17'd4658: data = 8'h02;
      17'd4659: data = 8'h2b;
      17'd4660: data = 8'hc5;
      17'd4661: data = 8'h06;
      17'd4662: data = 8'h33;
      17'd4663: data = 8'hcb;
      17'd4664: data = 8'h01;
      17'd4665: data = 8'h24;
      17'd4666: data = 8'hdb;
      17'd4667: data = 8'h06;
      17'd4668: data = 8'h0c;
      17'd4669: data = 8'hfd;
      17'd4670: data = 8'h02;
      17'd4671: data = 8'hd3;
      17'd4672: data = 8'h2d;
      17'd4673: data = 8'h16;
      17'd4674: data = 8'hc5;
      17'd4675: data = 8'h1f;
      17'd4676: data = 8'h01;
      17'd4677: data = 8'hdc;
      17'd4678: data = 8'h26;
      17'd4679: data = 8'hfd;
      17'd4680: data = 8'he2;
      17'd4681: data = 8'h1b;
      17'd4682: data = 8'h00;
      17'd4683: data = 8'hd5;
      17'd4684: data = 8'hfc;
      17'd4685: data = 8'h2d;
      17'd4686: data = 8'h00;
      17'd4687: data = 8'hce;
      17'd4688: data = 8'hfe;
      17'd4689: data = 8'h0e;
      17'd4690: data = 8'h1e;
      17'd4691: data = 8'hfc;
      17'd4692: data = 8'hce;
      17'd4693: data = 8'h1b;
      17'd4694: data = 8'h19;
      17'd4695: data = 8'he7;
      17'd4696: data = 8'hf2;
      17'd4697: data = 8'h0c;
      17'd4698: data = 8'h13;
      17'd4699: data = 8'heb;
      17'd4700: data = 8'hf2;
      17'd4701: data = 8'h13;
      17'd4702: data = 8'h0a;
      17'd4703: data = 8'h09;
      17'd4704: data = 8'heb;
      17'd4705: data = 8'h04;
      17'd4706: data = 8'h1b;
      17'd4707: data = 8'hd8;
      17'd4708: data = 8'h09;
      17'd4709: data = 8'h13;
      17'd4710: data = 8'hd8;
      17'd4711: data = 8'h09;
      17'd4712: data = 8'h0e;
      17'd4713: data = 8'hf6;
      17'd4714: data = 8'hfa;
      17'd4715: data = 8'h00;
      17'd4716: data = 8'h29;
      17'd4717: data = 8'hf9;
      17'd4718: data = 8'he7;
      17'd4719: data = 8'h13;
      17'd4720: data = 8'he5;
      17'd4721: data = 8'h11;
      17'd4722: data = 8'h22;
      17'd4723: data = 8'hd1;
      17'd4724: data = 8'hfe;
      17'd4725: data = 8'h11;
      17'd4726: data = 8'hec;
      17'd4727: data = 8'h16;
      17'd4728: data = 8'h1e;
      17'd4729: data = 8'he2;
      17'd4730: data = 8'he0;
      17'd4731: data = 8'h2c;
      17'd4732: data = 8'h0e;
      17'd4733: data = 8'hd8;
      17'd4734: data = 8'hfd;
      17'd4735: data = 8'h15;
      17'd4736: data = 8'hf2;
      17'd4737: data = 8'he7;
      17'd4738: data = 8'h1f;
      17'd4739: data = 8'h02;
      17'd4740: data = 8'hd8;
      17'd4741: data = 8'h1b;
      17'd4742: data = 8'h27;
      17'd4743: data = 8'he0;
      17'd4744: data = 8'he7;
      17'd4745: data = 8'h1f;
      17'd4746: data = 8'hfe;
      17'd4747: data = 8'h06;
      17'd4748: data = 8'h09;
      17'd4749: data = 8'hce;
      17'd4750: data = 8'h09;
      17'd4751: data = 8'h2d;
      17'd4752: data = 8'hf2;
      17'd4753: data = 8'hf1;
      17'd4754: data = 8'h02;
      17'd4755: data = 8'h01;
      17'd4756: data = 8'h0c;
      17'd4757: data = 8'h0d;
      17'd4758: data = 8'hfe;
      17'd4759: data = 8'he0;
      17'd4760: data = 8'h01;
      17'd4761: data = 8'h1c;
      17'd4762: data = 8'hed;
      17'd4763: data = 8'hf5;
      17'd4764: data = 8'h0d;
      17'd4765: data = 8'hfa;
      17'd4766: data = 8'hf6;
      17'd4767: data = 8'h13;
      17'd4768: data = 8'h01;
      17'd4769: data = 8'hf9;
      17'd4770: data = 8'h11;
      17'd4771: data = 8'hf2;
      17'd4772: data = 8'hfe;
      17'd4773: data = 8'h13;
      17'd4774: data = 8'hf4;
      17'd4775: data = 8'hef;
      17'd4776: data = 8'h0e;
      17'd4777: data = 8'h0e;
      17'd4778: data = 8'he5;
      17'd4779: data = 8'hec;
      17'd4780: data = 8'h16;
      17'd4781: data = 8'h12;
      17'd4782: data = 8'he9;
      17'd4783: data = 8'hfd;
      17'd4784: data = 8'h02;
      17'd4785: data = 8'hf6;
      17'd4786: data = 8'h06;
      17'd4787: data = 8'heb;
      17'd4788: data = 8'hfc;
      17'd4789: data = 8'h0e;
      17'd4790: data = 8'hf4;
      17'd4791: data = 8'hfa;
      17'd4792: data = 8'hf6;
      17'd4793: data = 8'h12;
      17'd4794: data = 8'h06;
      17'd4795: data = 8'heb;
      17'd4796: data = 8'hf6;
      17'd4797: data = 8'hf5;
      17'd4798: data = 8'h0e;
      17'd4799: data = 8'hfd;
      17'd4800: data = 8'hed;
      17'd4801: data = 8'h06;
      17'd4802: data = 8'hfd;
      17'd4803: data = 8'hf9;
      17'd4804: data = 8'hfa;
      17'd4805: data = 8'h1b;
      17'd4806: data = 8'h0d;
      17'd4807: data = 8'hd1;
      17'd4808: data = 8'h00;
      17'd4809: data = 8'h1f;
      17'd4810: data = 8'h09;
      17'd4811: data = 8'he7;
      17'd4812: data = 8'hf2;
      17'd4813: data = 8'h13;
      17'd4814: data = 8'hfa;
      17'd4815: data = 8'h09;
      17'd4816: data = 8'hf6;
      17'd4817: data = 8'he7;
      17'd4818: data = 8'h1e;
      17'd4819: data = 8'h0e;
      17'd4820: data = 8'he0;
      17'd4821: data = 8'h02;
      17'd4822: data = 8'h11;
      17'd4823: data = 8'hf5;
      17'd4824: data = 8'hfa;
      17'd4825: data = 8'h16;
      17'd4826: data = 8'h06;
      17'd4827: data = 8'hd6;
      17'd4828: data = 8'h05;
      17'd4829: data = 8'h1a;
      17'd4830: data = 8'h04;
      17'd4831: data = 8'hfd;
      17'd4832: data = 8'hf5;
      17'd4833: data = 8'hec;
      17'd4834: data = 8'h09;
      17'd4835: data = 8'h1e;
      17'd4836: data = 8'hf2;
      17'd4837: data = 8'he5;
      17'd4838: data = 8'h09;
      17'd4839: data = 8'h05;
      17'd4840: data = 8'hec;
      17'd4841: data = 8'h0d;
      17'd4842: data = 8'h13;
      17'd4843: data = 8'he3;
      17'd4844: data = 8'hf6;
      17'd4845: data = 8'h13;
      17'd4846: data = 8'hf1;
      17'd4847: data = 8'hf2;
      17'd4848: data = 8'h15;
      17'd4849: data = 8'h02;
      17'd4850: data = 8'heb;
      17'd4851: data = 8'h04;
      17'd4852: data = 8'h05;
      17'd4853: data = 8'h00;
      17'd4854: data = 8'h16;
      17'd4855: data = 8'h00;
      17'd4856: data = 8'hef;
      17'd4857: data = 8'hf6;
      17'd4858: data = 8'h04;
      17'd4859: data = 8'h0c;
      17'd4860: data = 8'hfa;
      17'd4861: data = 8'h00;
      17'd4862: data = 8'h00;
      17'd4863: data = 8'he9;
      17'd4864: data = 8'hfe;
      17'd4865: data = 8'h19;
      17'd4866: data = 8'h13;
      17'd4867: data = 8'hec;
      17'd4868: data = 8'hf4;
      17'd4869: data = 8'h15;
      17'd4870: data = 8'hfa;
      17'd4871: data = 8'hfd;
      17'd4872: data = 8'h04;
      17'd4873: data = 8'hf9;
      17'd4874: data = 8'hf6;
      17'd4875: data = 8'h01;
      17'd4876: data = 8'hf6;
      17'd4877: data = 8'h04;
      17'd4878: data = 8'h0c;
      17'd4879: data = 8'hfa;
      17'd4880: data = 8'h04;
      17'd4881: data = 8'hf6;
      17'd4882: data = 8'h01;
      17'd4883: data = 8'h0a;
      17'd4884: data = 8'hf5;
      17'd4885: data = 8'h00;
      17'd4886: data = 8'h01;
      17'd4887: data = 8'hef;
      17'd4888: data = 8'hf1;
      17'd4889: data = 8'h09;
      17'd4890: data = 8'h1c;
      17'd4891: data = 8'he9;
      17'd4892: data = 8'he7;
      17'd4893: data = 8'h1a;
      17'd4894: data = 8'h06;
      17'd4895: data = 8'he9;
      17'd4896: data = 8'hfc;
      17'd4897: data = 8'h15;
      17'd4898: data = 8'hfc;
      17'd4899: data = 8'he4;
      17'd4900: data = 8'hf5;
      17'd4901: data = 8'h0e;
      17'd4902: data = 8'h13;
      17'd4903: data = 8'hf4;
      17'd4904: data = 8'hf4;
      17'd4905: data = 8'h00;
      17'd4906: data = 8'hf6;
      17'd4907: data = 8'h15;
      17'd4908: data = 8'h0a;
      17'd4909: data = 8'hed;
      17'd4910: data = 8'hfc;
      17'd4911: data = 8'h0e;
      17'd4912: data = 8'hfe;
      17'd4913: data = 8'hfe;
      17'd4914: data = 8'h11;
      17'd4915: data = 8'hf9;
      17'd4916: data = 8'hfa;
      17'd4917: data = 8'h09;
      17'd4918: data = 8'h02;
      17'd4919: data = 8'hfa;
      17'd4920: data = 8'hfd;
      17'd4921: data = 8'h11;
      17'd4922: data = 8'h05;
      17'd4923: data = 8'he5;
      17'd4924: data = 8'h01;
      17'd4925: data = 8'h0c;
      17'd4926: data = 8'hf4;
      17'd4927: data = 8'h05;
      17'd4928: data = 8'h0d;
      17'd4929: data = 8'hf5;
      17'd4930: data = 8'hf2;
      17'd4931: data = 8'h15;
      17'd4932: data = 8'h06;
      17'd4933: data = 8'hed;
      17'd4934: data = 8'hfe;
      17'd4935: data = 8'h05;
      17'd4936: data = 8'h02;
      17'd4937: data = 8'h02;
      17'd4938: data = 8'hf9;
      17'd4939: data = 8'h09;
      17'd4940: data = 8'h0c;
      17'd4941: data = 8'hf6;
      17'd4942: data = 8'h02;
      17'd4943: data = 8'h00;
      17'd4944: data = 8'hfa;
      17'd4945: data = 8'hfe;
      17'd4946: data = 8'h0e;
      17'd4947: data = 8'h00;
      17'd4948: data = 8'heb;
      17'd4949: data = 8'hfe;
      17'd4950: data = 8'h06;
      17'd4951: data = 8'h04;
      17'd4952: data = 8'h0c;
      17'd4953: data = 8'hf9;
      17'd4954: data = 8'hef;
      17'd4955: data = 8'h1c;
      17'd4956: data = 8'h09;
      17'd4957: data = 8'hf1;
      17'd4958: data = 8'h04;
      17'd4959: data = 8'hf9;
      17'd4960: data = 8'hf9;
      17'd4961: data = 8'hfe;
      17'd4962: data = 8'h00;
      17'd4963: data = 8'h06;
      17'd4964: data = 8'hf4;
      17'd4965: data = 8'h12;
      17'd4966: data = 8'h09;
      17'd4967: data = 8'he2;
      17'd4968: data = 8'h0c;
      17'd4969: data = 8'h11;
      17'd4970: data = 8'hf5;
      17'd4971: data = 8'hfc;
      17'd4972: data = 8'h0d;
      17'd4973: data = 8'hf9;
      17'd4974: data = 8'hfa;
      17'd4975: data = 8'h11;
      17'd4976: data = 8'h02;
      17'd4977: data = 8'heb;
      17'd4978: data = 8'h05;
      17'd4979: data = 8'h0c;
      17'd4980: data = 8'hf5;
      17'd4981: data = 8'h11;
      17'd4982: data = 8'h04;
      17'd4983: data = 8'hec;
      17'd4984: data = 8'h04;
      17'd4985: data = 8'h16;
      17'd4986: data = 8'hed;
      17'd4987: data = 8'hf1;
      17'd4988: data = 8'h13;
      17'd4989: data = 8'hfd;
      17'd4990: data = 8'hec;
      17'd4991: data = 8'h01;
      17'd4992: data = 8'h0a;
      17'd4993: data = 8'h00;
      17'd4994: data = 8'hfe;
      17'd4995: data = 8'hfd;
      17'd4996: data = 8'hed;
      17'd4997: data = 8'hf2;
      17'd4998: data = 8'h06;
      17'd4999: data = 8'h04;
      17'd5000: data = 8'h01;
      17'd5001: data = 8'hfc;
      17'd5002: data = 8'hf2;
      17'd5003: data = 8'hf5;
      17'd5004: data = 8'h04;
      17'd5005: data = 8'h0d;
      17'd5006: data = 8'hf9;
      17'd5007: data = 8'hf5;
      17'd5008: data = 8'hf6;
      17'd5009: data = 8'hfc;
      17'd5010: data = 8'h09;
      17'd5011: data = 8'h02;
      17'd5012: data = 8'hef;
      17'd5013: data = 8'hfa;
      17'd5014: data = 8'h06;
      17'd5015: data = 8'hfa;
      17'd5016: data = 8'h00;
      17'd5017: data = 8'h06;
      17'd5018: data = 8'h01;
      17'd5019: data = 8'hf6;
      17'd5020: data = 8'hfd;
      17'd5021: data = 8'hfd;
      17'd5022: data = 8'hf6;
      17'd5023: data = 8'h00;
      17'd5024: data = 8'h05;
      17'd5025: data = 8'h02;
      17'd5026: data = 8'hf5;
      17'd5027: data = 8'hfa;
      17'd5028: data = 8'h02;
      17'd5029: data = 8'h02;
      17'd5030: data = 8'h00;
      17'd5031: data = 8'hfe;
      17'd5032: data = 8'hfa;
      17'd5033: data = 8'hf5;
      17'd5034: data = 8'h04;
      17'd5035: data = 8'h11;
      17'd5036: data = 8'hfe;
      17'd5037: data = 8'hf6;
      17'd5038: data = 8'hfa;
      17'd5039: data = 8'hfe;
      17'd5040: data = 8'h0d;
      17'd5041: data = 8'h02;
      17'd5042: data = 8'hf6;
      17'd5043: data = 8'hfc;
      17'd5044: data = 8'h09;
      17'd5045: data = 8'h04;
      17'd5046: data = 8'hf6;
      17'd5047: data = 8'hf6;
      17'd5048: data = 8'hfe;
      17'd5049: data = 8'h06;
      17'd5050: data = 8'hfa;
      17'd5051: data = 8'hf6;
      17'd5052: data = 8'h06;
      17'd5053: data = 8'h04;
      17'd5054: data = 8'h00;
      17'd5055: data = 8'h00;
      17'd5056: data = 8'hf6;
      17'd5057: data = 8'hf4;
      17'd5058: data = 8'hf4;
      17'd5059: data = 8'h01;
      17'd5060: data = 8'h06;
      17'd5061: data = 8'hfc;
      17'd5062: data = 8'hfe;
      17'd5063: data = 8'hf9;
      17'd5064: data = 8'h04;
      17'd5065: data = 8'h06;
      17'd5066: data = 8'hf4;
      17'd5067: data = 8'hfa;
      17'd5068: data = 8'h09;
      17'd5069: data = 8'h05;
      17'd5070: data = 8'hf1;
      17'd5071: data = 8'hfa;
      17'd5072: data = 8'h06;
      17'd5073: data = 8'h01;
      17'd5074: data = 8'hfa;
      17'd5075: data = 8'hfc;
      17'd5076: data = 8'hfd;
      17'd5077: data = 8'hf9;
      17'd5078: data = 8'hfe;
      17'd5079: data = 8'h15;
      17'd5080: data = 8'h09;
      17'd5081: data = 8'hec;
      17'd5082: data = 8'hfc;
      17'd5083: data = 8'h02;
      17'd5084: data = 8'hfd;
      17'd5085: data = 8'hf9;
      17'd5086: data = 8'h01;
      17'd5087: data = 8'h01;
      17'd5088: data = 8'hf9;
      17'd5089: data = 8'h02;
      17'd5090: data = 8'h02;
      17'd5091: data = 8'h05;
      17'd5092: data = 8'h00;
      17'd5093: data = 8'hf2;
      17'd5094: data = 8'hfa;
      17'd5095: data = 8'h01;
      17'd5096: data = 8'h01;
      17'd5097: data = 8'hfc;
      17'd5098: data = 8'h01;
      17'd5099: data = 8'hfd;
      17'd5100: data = 8'hf9;
      17'd5101: data = 8'hfc;
      17'd5102: data = 8'hfd;
      17'd5103: data = 8'h00;
      17'd5104: data = 8'hfe;
      17'd5105: data = 8'h04;
      17'd5106: data = 8'h02;
      17'd5107: data = 8'h01;
      17'd5108: data = 8'hf9;
      17'd5109: data = 8'hfe;
      17'd5110: data = 8'h04;
      17'd5111: data = 8'hf9;
      17'd5112: data = 8'hf1;
      17'd5113: data = 8'hfc;
      17'd5114: data = 8'h0c;
      17'd5115: data = 8'h01;
      17'd5116: data = 8'hf6;
      17'd5117: data = 8'h05;
      17'd5118: data = 8'h02;
      17'd5119: data = 8'hf5;
      17'd5120: data = 8'hfe;
      17'd5121: data = 8'h02;
      17'd5122: data = 8'hfc;
      17'd5123: data = 8'hf6;
      17'd5124: data = 8'h0a;
      17'd5125: data = 8'h0a;
      17'd5126: data = 8'hf2;
      17'd5127: data = 8'hfd;
      17'd5128: data = 8'h01;
      17'd5129: data = 8'hfe;
      17'd5130: data = 8'h01;
      17'd5131: data = 8'hf9;
      17'd5132: data = 8'hf4;
      17'd5133: data = 8'h09;
      17'd5134: data = 8'h15;
      17'd5135: data = 8'hfe;
      17'd5136: data = 8'hf1;
      17'd5137: data = 8'hf6;
      17'd5138: data = 8'h05;
      17'd5139: data = 8'h06;
      17'd5140: data = 8'hfd;
      17'd5141: data = 8'hf4;
      17'd5142: data = 8'hfc;
      17'd5143: data = 8'h09;
      17'd5144: data = 8'h06;
      17'd5145: data = 8'hf9;
      17'd5146: data = 8'hf5;
      17'd5147: data = 8'h02;
      17'd5148: data = 8'hfe;
      17'd5149: data = 8'hfd;
      17'd5150: data = 8'h00;
      17'd5151: data = 8'hfe;
      17'd5152: data = 8'hfa;
      17'd5153: data = 8'h0a;
      17'd5154: data = 8'h11;
      17'd5155: data = 8'hf2;
      17'd5156: data = 8'hf4;
      17'd5157: data = 8'h01;
      17'd5158: data = 8'hfe;
      17'd5159: data = 8'h01;
      17'd5160: data = 8'hfd;
      17'd5161: data = 8'hfc;
      17'd5162: data = 8'h09;
      17'd5163: data = 8'h06;
      17'd5164: data = 8'h00;
      17'd5165: data = 8'h00;
      17'd5166: data = 8'h05;
      17'd5167: data = 8'hfc;
      17'd5168: data = 8'hf6;
      17'd5169: data = 8'h05;
      17'd5170: data = 8'h06;
      17'd5171: data = 8'hfd;
      17'd5172: data = 8'h02;
      17'd5173: data = 8'h0d;
      17'd5174: data = 8'hf9;
      17'd5175: data = 8'hf4;
      17'd5176: data = 8'h11;
      17'd5177: data = 8'h06;
      17'd5178: data = 8'hf9;
      17'd5179: data = 8'hfd;
      17'd5180: data = 8'hf9;
      17'd5181: data = 8'h06;
      17'd5182: data = 8'h0d;
      17'd5183: data = 8'h00;
      17'd5184: data = 8'hf6;
      17'd5185: data = 8'hef;
      17'd5186: data = 8'h05;
      17'd5187: data = 8'h0a;
      17'd5188: data = 8'hfe;
      17'd5189: data = 8'h01;
      17'd5190: data = 8'h06;
      17'd5191: data = 8'h0e;
      17'd5192: data = 8'h00;
      17'd5193: data = 8'hfc;
      17'd5194: data = 8'h02;
      17'd5195: data = 8'hf9;
      17'd5196: data = 8'h01;
      17'd5197: data = 8'h09;
      17'd5198: data = 8'hfe;
      17'd5199: data = 8'hf9;
      17'd5200: data = 8'h06;
      17'd5201: data = 8'h0d;
      17'd5202: data = 8'h01;
      17'd5203: data = 8'hfc;
      17'd5204: data = 8'hf5;
      17'd5205: data = 8'hfd;
      17'd5206: data = 8'h0e;
      17'd5207: data = 8'h00;
      17'd5208: data = 8'hf2;
      17'd5209: data = 8'h02;
      17'd5210: data = 8'h00;
      17'd5211: data = 8'hfe;
      17'd5212: data = 8'hfd;
      17'd5213: data = 8'hf6;
      17'd5214: data = 8'hfd;
      17'd5215: data = 8'hfe;
      17'd5216: data = 8'h01;
      17'd5217: data = 8'h05;
      17'd5218: data = 8'hfe;
      17'd5219: data = 8'hfa;
      17'd5220: data = 8'h00;
      17'd5221: data = 8'hfe;
      17'd5222: data = 8'hfc;
      17'd5223: data = 8'hf9;
      17'd5224: data = 8'hfd;
      17'd5225: data = 8'h00;
      17'd5226: data = 8'h01;
      17'd5227: data = 8'h02;
      17'd5228: data = 8'hfe;
      17'd5229: data = 8'h00;
      17'd5230: data = 8'h00;
      17'd5231: data = 8'hfe;
      17'd5232: data = 8'h02;
      17'd5233: data = 8'h01;
      17'd5234: data = 8'hfc;
      17'd5235: data = 8'hfd;
      17'd5236: data = 8'h00;
      17'd5237: data = 8'h01;
      17'd5238: data = 8'h04;
      17'd5239: data = 8'h01;
      17'd5240: data = 8'hfd;
      17'd5241: data = 8'hfe;
      17'd5242: data = 8'h00;
      17'd5243: data = 8'h02;
      17'd5244: data = 8'h04;
      17'd5245: data = 8'h05;
      17'd5246: data = 8'h02;
      17'd5247: data = 8'hfe;
      17'd5248: data = 8'hfe;
      17'd5249: data = 8'h01;
      17'd5250: data = 8'h04;
      17'd5251: data = 8'h00;
      17'd5252: data = 8'hfe;
      17'd5253: data = 8'h00;
      17'd5254: data = 8'h06;
      17'd5255: data = 8'h05;
      17'd5256: data = 8'h01;
      17'd5257: data = 8'h01;
      17'd5258: data = 8'h00;
      17'd5259: data = 8'h01;
      17'd5260: data = 8'hfc;
      17'd5261: data = 8'hfe;
      17'd5262: data = 8'h05;
      17'd5263: data = 8'h01;
      17'd5264: data = 8'h01;
      17'd5265: data = 8'hfe;
      17'd5266: data = 8'hfe;
      17'd5267: data = 8'h00;
      17'd5268: data = 8'hfe;
      17'd5269: data = 8'hfe;
      17'd5270: data = 8'hfc;
      17'd5271: data = 8'hfe;
      17'd5272: data = 8'h00;
      17'd5273: data = 8'hfd;
      17'd5274: data = 8'h04;
      17'd5275: data = 8'h02;
      17'd5276: data = 8'hfc;
      17'd5277: data = 8'hfe;
      17'd5278: data = 8'h00;
      17'd5279: data = 8'h00;
      17'd5280: data = 8'h04;
      17'd5281: data = 8'h01;
      17'd5282: data = 8'hf9;
      17'd5283: data = 8'hfc;
      17'd5284: data = 8'h00;
      17'd5285: data = 8'h00;
      17'd5286: data = 8'hf9;
      17'd5287: data = 8'hfd;
      17'd5288: data = 8'h04;
      17'd5289: data = 8'hfd;
      17'd5290: data = 8'hfd;
      17'd5291: data = 8'h02;
      17'd5292: data = 8'h02;
      17'd5293: data = 8'hfe;
      17'd5294: data = 8'h01;
      17'd5295: data = 8'h00;
      17'd5296: data = 8'hfc;
      17'd5297: data = 8'hfa;
      17'd5298: data = 8'hfe;
      17'd5299: data = 8'h02;
      17'd5300: data = 8'h00;
      17'd5301: data = 8'hfa;
      17'd5302: data = 8'hfe;
      17'd5303: data = 8'h04;
      17'd5304: data = 8'hfe;
      17'd5305: data = 8'hfc;
      17'd5306: data = 8'hf6;
      17'd5307: data = 8'hf6;
      17'd5308: data = 8'hfc;
      17'd5309: data = 8'hfd;
      17'd5310: data = 8'h00;
      17'd5311: data = 8'hf1;
      17'd5312: data = 8'hf1;
      17'd5313: data = 8'hf6;
      17'd5314: data = 8'hf9;
      17'd5315: data = 8'hfa;
      17'd5316: data = 8'hf4;
      17'd5317: data = 8'h00;
      17'd5318: data = 8'h00;
      17'd5319: data = 8'hf4;
      17'd5320: data = 8'hf6;
      17'd5321: data = 8'hfc;
      17'd5322: data = 8'hf5;
      17'd5323: data = 8'hf6;
      17'd5324: data = 8'h01;
      17'd5325: data = 8'hfc;
      17'd5326: data = 8'hf6;
      17'd5327: data = 8'h04;
      17'd5328: data = 8'h04;
      17'd5329: data = 8'h05;
      17'd5330: data = 8'h11;
      17'd5331: data = 8'h02;
      17'd5332: data = 8'hfc;
      17'd5333: data = 8'h05;
      17'd5334: data = 8'h0d;
      17'd5335: data = 8'h09;
      17'd5336: data = 8'h04;
      17'd5337: data = 8'h0d;
      17'd5338: data = 8'h04;
      17'd5339: data = 8'h04;
      17'd5340: data = 8'h0d;
      17'd5341: data = 8'h09;
      17'd5342: data = 8'h0d;
      17'd5343: data = 8'h11;
      17'd5344: data = 8'h0c;
      17'd5345: data = 8'h0a;
      17'd5346: data = 8'h06;
      17'd5347: data = 8'h05;
      17'd5348: data = 8'h0c;
      17'd5349: data = 8'h0c;
      17'd5350: data = 8'h06;
      17'd5351: data = 8'h06;
      17'd5352: data = 8'h02;
      17'd5353: data = 8'hfc;
      17'd5354: data = 8'h04;
      17'd5355: data = 8'h12;
      17'd5356: data = 8'h05;
      17'd5357: data = 8'hfe;
      17'd5358: data = 8'hf9;
      17'd5359: data = 8'h00;
      17'd5360: data = 8'h09;
      17'd5361: data = 8'h06;
      17'd5362: data = 8'h00;
      17'd5363: data = 8'hf9;
      17'd5364: data = 8'hf9;
      17'd5365: data = 8'hf4;
      17'd5366: data = 8'h01;
      17'd5367: data = 8'h00;
      17'd5368: data = 8'hf1;
      17'd5369: data = 8'hf1;
      17'd5370: data = 8'hf9;
      17'd5371: data = 8'hf6;
      17'd5372: data = 8'hfc;
      17'd5373: data = 8'hf6;
      17'd5374: data = 8'hed;
      17'd5375: data = 8'hf6;
      17'd5376: data = 8'hf5;
      17'd5377: data = 8'hfc;
      17'd5378: data = 8'hf2;
      17'd5379: data = 8'hf1;
      17'd5380: data = 8'hf2;
      17'd5381: data = 8'hf5;
      17'd5382: data = 8'h04;
      17'd5383: data = 8'hf5;
      17'd5384: data = 8'hec;
      17'd5385: data = 8'hf4;
      17'd5386: data = 8'hf9;
      17'd5387: data = 8'hfd;
      17'd5388: data = 8'hfc;
      17'd5389: data = 8'hec;
      17'd5390: data = 8'hf1;
      17'd5391: data = 8'hfc;
      17'd5392: data = 8'hf6;
      17'd5393: data = 8'hfa;
      17'd5394: data = 8'hfa;
      17'd5395: data = 8'hf4;
      17'd5396: data = 8'hfd;
      17'd5397: data = 8'h0a;
      17'd5398: data = 8'h02;
      17'd5399: data = 8'hf4;
      17'd5400: data = 8'hf6;
      17'd5401: data = 8'hf6;
      17'd5402: data = 8'hef;
      17'd5403: data = 8'hf2;
      17'd5404: data = 8'hfa;
      17'd5405: data = 8'hf9;
      17'd5406: data = 8'h05;
      17'd5407: data = 8'h11;
      17'd5408: data = 8'h02;
      17'd5409: data = 8'hfd;
      17'd5410: data = 8'hfe;
      17'd5411: data = 8'hfe;
      17'd5412: data = 8'hfa;
      17'd5413: data = 8'hfc;
      17'd5414: data = 8'hf9;
      17'd5415: data = 8'hfc;
      17'd5416: data = 8'h06;
      17'd5417: data = 8'h05;
      17'd5418: data = 8'hfe;
      17'd5419: data = 8'h05;
      17'd5420: data = 8'h05;
      17'd5421: data = 8'h01;
      17'd5422: data = 8'h0a;
      17'd5423: data = 8'h06;
      17'd5424: data = 8'h01;
      17'd5425: data = 8'h05;
      17'd5426: data = 8'h0a;
      17'd5427: data = 8'h04;
      17'd5428: data = 8'h01;
      17'd5429: data = 8'h06;
      17'd5430: data = 8'h09;
      17'd5431: data = 8'h09;
      17'd5432: data = 8'h12;
      17'd5433: data = 8'h0e;
      17'd5434: data = 8'h09;
      17'd5435: data = 8'h11;
      17'd5436: data = 8'h0a;
      17'd5437: data = 8'h02;
      17'd5438: data = 8'h01;
      17'd5439: data = 8'h00;
      17'd5440: data = 8'hfe;
      17'd5441: data = 8'h06;
      17'd5442: data = 8'h0e;
      17'd5443: data = 8'h0e;
      17'd5444: data = 8'h0c;
      17'd5445: data = 8'h02;
      17'd5446: data = 8'h04;
      17'd5447: data = 8'h02;
      17'd5448: data = 8'hfc;
      17'd5449: data = 8'hfc;
      17'd5450: data = 8'hfa;
      17'd5451: data = 8'hfa;
      17'd5452: data = 8'hfc;
      17'd5453: data = 8'hf6;
      17'd5454: data = 8'hfd;
      17'd5455: data = 8'hfe;
      17'd5456: data = 8'hfc;
      17'd5457: data = 8'hf9;
      17'd5458: data = 8'hf9;
      17'd5459: data = 8'hfd;
      17'd5460: data = 8'hfe;
      17'd5461: data = 8'hf6;
      17'd5462: data = 8'hef;
      17'd5463: data = 8'hf1;
      17'd5464: data = 8'hef;
      17'd5465: data = 8'hec;
      17'd5466: data = 8'hec;
      17'd5467: data = 8'hf4;
      17'd5468: data = 8'hfe;
      17'd5469: data = 8'hf5;
      17'd5470: data = 8'hed;
      17'd5471: data = 8'hfa;
      17'd5472: data = 8'hf6;
      17'd5473: data = 8'hed;
      17'd5474: data = 8'hed;
      17'd5475: data = 8'hed;
      17'd5476: data = 8'hf1;
      17'd5477: data = 8'hf9;
      17'd5478: data = 8'hf9;
      17'd5479: data = 8'hfd;
      17'd5480: data = 8'h04;
      17'd5481: data = 8'h01;
      17'd5482: data = 8'hfd;
      17'd5483: data = 8'h04;
      17'd5484: data = 8'h09;
      17'd5485: data = 8'h00;
      17'd5486: data = 8'h04;
      17'd5487: data = 8'h15;
      17'd5488: data = 8'h15;
      17'd5489: data = 8'h11;
      17'd5490: data = 8'h23;
      17'd5491: data = 8'h27;
      17'd5492: data = 8'h1a;
      17'd5493: data = 8'h1b;
      17'd5494: data = 8'h27;
      17'd5495: data = 8'h1f;
      17'd5496: data = 8'h23;
      17'd5497: data = 8'h24;
      17'd5498: data = 8'h1f;
      17'd5499: data = 8'h23;
      17'd5500: data = 8'h26;
      17'd5501: data = 8'h27;
      17'd5502: data = 8'h27;
      17'd5503: data = 8'h27;
      17'd5504: data = 8'h29;
      17'd5505: data = 8'h22;
      17'd5506: data = 8'h22;
      17'd5507: data = 8'h1f;
      17'd5508: data = 8'h1b;
      17'd5509: data = 8'h1a;
      17'd5510: data = 8'h13;
      17'd5511: data = 8'h16;
      17'd5512: data = 8'h12;
      17'd5513: data = 8'h0d;
      17'd5514: data = 8'h12;
      17'd5515: data = 8'h13;
      17'd5516: data = 8'h0d;
      17'd5517: data = 8'h02;
      17'd5518: data = 8'h02;
      17'd5519: data = 8'h01;
      17'd5520: data = 8'hf9;
      17'd5521: data = 8'hfa;
      17'd5522: data = 8'hf2;
      17'd5523: data = 8'hf2;
      17'd5524: data = 8'hf5;
      17'd5525: data = 8'he4;
      17'd5526: data = 8'heb;
      17'd5527: data = 8'hf6;
      17'd5528: data = 8'he7;
      17'd5529: data = 8'hda;
      17'd5530: data = 8'hde;
      17'd5531: data = 8'he0;
      17'd5532: data = 8'hd5;
      17'd5533: data = 8'hd5;
      17'd5534: data = 8'hd1;
      17'd5535: data = 8'hd2;
      17'd5536: data = 8'hd3;
      17'd5537: data = 8'hc6;
      17'd5538: data = 8'hd2;
      17'd5539: data = 8'he9;
      17'd5540: data = 8'he0;
      17'd5541: data = 8'hd8;
      17'd5542: data = 8'hc4;
      17'd5543: data = 8'hc6;
      17'd5544: data = 8'he2;
      17'd5545: data = 8'hc6;
      17'd5546: data = 8'hd3;
      17'd5547: data = 8'he4;
      17'd5548: data = 8'he3;
      17'd5549: data = 8'heb;
      17'd5550: data = 8'hde;
      17'd5551: data = 8'he9;
      17'd5552: data = 8'heb;
      17'd5553: data = 8'hed;
      17'd5554: data = 8'hfd;
      17'd5555: data = 8'hf1;
      17'd5556: data = 8'hf5;
      17'd5557: data = 8'h00;
      17'd5558: data = 8'hfa;
      17'd5559: data = 8'h04;
      17'd5560: data = 8'h09;
      17'd5561: data = 8'h00;
      17'd5562: data = 8'hf5;
      17'd5563: data = 8'h01;
      17'd5564: data = 8'h13;
      17'd5565: data = 8'h13;
      17'd5566: data = 8'h12;
      17'd5567: data = 8'h12;
      17'd5568: data = 8'h13;
      17'd5569: data = 8'h05;
      17'd5570: data = 8'h09;
      17'd5571: data = 8'h0d;
      17'd5572: data = 8'h04;
      17'd5573: data = 8'h13;
      17'd5574: data = 8'h0e;
      17'd5575: data = 8'h0d;
      17'd5576: data = 8'h16;
      17'd5577: data = 8'h11;
      17'd5578: data = 8'h0e;
      17'd5579: data = 8'h0c;
      17'd5580: data = 8'h04;
      17'd5581: data = 8'hf6;
      17'd5582: data = 8'hf9;
      17'd5583: data = 8'h09;
      17'd5584: data = 8'h0d;
      17'd5585: data = 8'h0c;
      17'd5586: data = 8'h00;
      17'd5587: data = 8'hf5;
      17'd5588: data = 8'h01;
      17'd5589: data = 8'h05;
      17'd5590: data = 8'hf9;
      17'd5591: data = 8'hf4;
      17'd5592: data = 8'hfa;
      17'd5593: data = 8'hf2;
      17'd5594: data = 8'he0;
      17'd5595: data = 8'hf1;
      17'd5596: data = 8'hf5;
      17'd5597: data = 8'he7;
      17'd5598: data = 8'hed;
      17'd5599: data = 8'hf4;
      17'd5600: data = 8'hec;
      17'd5601: data = 8'hec;
      17'd5602: data = 8'hf2;
      17'd5603: data = 8'hf1;
      17'd5604: data = 8'hfa;
      17'd5605: data = 8'hfc;
      17'd5606: data = 8'hed;
      17'd5607: data = 8'hec;
      17'd5608: data = 8'hf2;
      17'd5609: data = 8'hf5;
      17'd5610: data = 8'hf9;
      17'd5611: data = 8'hf5;
      17'd5612: data = 8'hfd;
      17'd5613: data = 8'h13;
      17'd5614: data = 8'h11;
      17'd5615: data = 8'hfc;
      17'd5616: data = 8'h05;
      17'd5617: data = 8'h0a;
      17'd5618: data = 8'h00;
      17'd5619: data = 8'h02;
      17'd5620: data = 8'h0c;
      17'd5621: data = 8'h11;
      17'd5622: data = 8'h13;
      17'd5623: data = 8'h1a;
      17'd5624: data = 8'h15;
      17'd5625: data = 8'h12;
      17'd5626: data = 8'h16;
      17'd5627: data = 8'h1c;
      17'd5628: data = 8'h1f;
      17'd5629: data = 8'h1b;
      17'd5630: data = 8'h16;
      17'd5631: data = 8'h15;
      17'd5632: data = 8'h12;
      17'd5633: data = 8'h16;
      17'd5634: data = 8'h1c;
      17'd5635: data = 8'h1a;
      17'd5636: data = 8'h13;
      17'd5637: data = 8'h12;
      17'd5638: data = 8'h19;
      17'd5639: data = 8'h1e;
      17'd5640: data = 8'h16;
      17'd5641: data = 8'h13;
      17'd5642: data = 8'h0e;
      17'd5643: data = 8'h04;
      17'd5644: data = 8'h02;
      17'd5645: data = 8'h01;
      17'd5646: data = 8'h00;
      17'd5647: data = 8'h00;
      17'd5648: data = 8'h04;
      17'd5649: data = 8'hfe;
      17'd5650: data = 8'hfd;
      17'd5651: data = 8'hfd;
      17'd5652: data = 8'hf6;
      17'd5653: data = 8'hf2;
      17'd5654: data = 8'hf1;
      17'd5655: data = 8'hf2;
      17'd5656: data = 8'hec;
      17'd5657: data = 8'he9;
      17'd5658: data = 8'hef;
      17'd5659: data = 8'hf2;
      17'd5660: data = 8'he9;
      17'd5661: data = 8'he4;
      17'd5662: data = 8'hec;
      17'd5663: data = 8'hef;
      17'd5664: data = 8'hf4;
      17'd5665: data = 8'hf1;
      17'd5666: data = 8'hed;
      17'd5667: data = 8'hf2;
      17'd5668: data = 8'hf5;
      17'd5669: data = 8'hf2;
      17'd5670: data = 8'hf1;
      17'd5671: data = 8'hf9;
      17'd5672: data = 8'h00;
      17'd5673: data = 8'hfe;
      17'd5674: data = 8'hfe;
      17'd5675: data = 8'h06;
      17'd5676: data = 8'h0d;
      17'd5677: data = 8'h0c;
      17'd5678: data = 8'h0c;
      17'd5679: data = 8'h0a;
      17'd5680: data = 8'h0c;
      17'd5681: data = 8'h12;
      17'd5682: data = 8'h12;
      17'd5683: data = 8'h1b;
      17'd5684: data = 8'h1f;
      17'd5685: data = 8'h1b;
      17'd5686: data = 8'h23;
      17'd5687: data = 8'h22;
      17'd5688: data = 8'h1a;
      17'd5689: data = 8'h23;
      17'd5690: data = 8'h24;
      17'd5691: data = 8'h1b;
      17'd5692: data = 8'h1e;
      17'd5693: data = 8'h24;
      17'd5694: data = 8'h23;
      17'd5695: data = 8'h26;
      17'd5696: data = 8'h29;
      17'd5697: data = 8'h29;
      17'd5698: data = 8'h2b;
      17'd5699: data = 8'h24;
      17'd5700: data = 8'h1c;
      17'd5701: data = 8'h1c;
      17'd5702: data = 8'h1c;
      17'd5703: data = 8'h1a;
      17'd5704: data = 8'h1a;
      17'd5705: data = 8'h1a;
      17'd5706: data = 8'h1c;
      17'd5707: data = 8'h1c;
      17'd5708: data = 8'h1b;
      17'd5709: data = 8'h19;
      17'd5710: data = 8'h13;
      17'd5711: data = 8'h12;
      17'd5712: data = 8'h0a;
      17'd5713: data = 8'h0c;
      17'd5714: data = 8'h0c;
      17'd5715: data = 8'h01;
      17'd5716: data = 8'hfe;
      17'd5717: data = 8'h00;
      17'd5718: data = 8'hfe;
      17'd5719: data = 8'h00;
      17'd5720: data = 8'hfd;
      17'd5721: data = 8'hfa;
      17'd5722: data = 8'hfa;
      17'd5723: data = 8'hf4;
      17'd5724: data = 8'hf1;
      17'd5725: data = 8'heb;
      17'd5726: data = 8'hec;
      17'd5727: data = 8'he9;
      17'd5728: data = 8'hdb;
      17'd5729: data = 8'he0;
      17'd5730: data = 8'he4;
      17'd5731: data = 8'he0;
      17'd5732: data = 8'hdc;
      17'd5733: data = 8'he0;
      17'd5734: data = 8'hdb;
      17'd5735: data = 8'hd5;
      17'd5736: data = 8'hd1;
      17'd5737: data = 8'hd1;
      17'd5738: data = 8'hce;
      17'd5739: data = 8'hcb;
      17'd5740: data = 8'hca;
      17'd5741: data = 8'hca;
      17'd5742: data = 8'hd1;
      17'd5743: data = 8'hd2;
      17'd5744: data = 8'hc6;
      17'd5745: data = 8'hc4;
      17'd5746: data = 8'hca;
      17'd5747: data = 8'hca;
      17'd5748: data = 8'hc9;
      17'd5749: data = 8'hc6;
      17'd5750: data = 8'hc4;
      17'd5751: data = 8'hca;
      17'd5752: data = 8'hd2;
      17'd5753: data = 8'hd3;
      17'd5754: data = 8'hd2;
      17'd5755: data = 8'hca;
      17'd5756: data = 8'hda;
      17'd5757: data = 8'hf1;
      17'd5758: data = 8'he3;
      17'd5759: data = 8'hce;
      17'd5760: data = 8'hdc;
      17'd5761: data = 8'he3;
      17'd5762: data = 8'hdb;
      17'd5763: data = 8'hec;
      17'd5764: data = 8'hfe;
      17'd5765: data = 8'hf5;
      17'd5766: data = 8'hf1;
      17'd5767: data = 8'hfd;
      17'd5768: data = 8'hfc;
      17'd5769: data = 8'hfe;
      17'd5770: data = 8'h06;
      17'd5771: data = 8'hf9;
      17'd5772: data = 8'h00;
      17'd5773: data = 8'h09;
      17'd5774: data = 8'h04;
      17'd5775: data = 8'h05;
      17'd5776: data = 8'h0d;
      17'd5777: data = 8'h0e;
      17'd5778: data = 8'h05;
      17'd5779: data = 8'h13;
      17'd5780: data = 8'h12;
      17'd5781: data = 8'h15;
      17'd5782: data = 8'h15;
      17'd5783: data = 8'h09;
      17'd5784: data = 8'h1a;
      17'd5785: data = 8'h12;
      17'd5786: data = 8'h05;
      17'd5787: data = 8'h09;
      17'd5788: data = 8'h19;
      17'd5789: data = 8'h11;
      17'd5790: data = 8'h16;
      17'd5791: data = 8'h15;
      17'd5792: data = 8'h01;
      17'd5793: data = 8'h05;
      17'd5794: data = 8'h0c;
      17'd5795: data = 8'h05;
      17'd5796: data = 8'h04;
      17'd5797: data = 8'h16;
      17'd5798: data = 8'h02;
      17'd5799: data = 8'hec;
      17'd5800: data = 8'hfd;
      17'd5801: data = 8'h00;
      17'd5802: data = 8'hf4;
      17'd5803: data = 8'hf2;
      17'd5804: data = 8'hf9;
      17'd5805: data = 8'hfe;
      17'd5806: data = 8'h00;
      17'd5807: data = 8'hfa;
      17'd5808: data = 8'hf1;
      17'd5809: data = 8'hed;
      17'd5810: data = 8'hfa;
      17'd5811: data = 8'hfe;
      17'd5812: data = 8'hf1;
      17'd5813: data = 8'hf5;
      17'd5814: data = 8'hfe;
      17'd5815: data = 8'hfc;
      17'd5816: data = 8'hf9;
      17'd5817: data = 8'hfc;
      17'd5818: data = 8'h00;
      17'd5819: data = 8'h01;
      17'd5820: data = 8'h0a;
      17'd5821: data = 8'h06;
      17'd5822: data = 8'h09;
      17'd5823: data = 8'h05;
      17'd5824: data = 8'hfe;
      17'd5825: data = 8'h0e;
      17'd5826: data = 8'h12;
      17'd5827: data = 8'h13;
      17'd5828: data = 8'h12;
      17'd5829: data = 8'h0d;
      17'd5830: data = 8'h16;
      17'd5831: data = 8'h13;
      17'd5832: data = 8'h15;
      17'd5833: data = 8'h1f;
      17'd5834: data = 8'h1e;
      17'd5835: data = 8'h1b;
      17'd5836: data = 8'h22;
      17'd5837: data = 8'h19;
      17'd5838: data = 8'h12;
      17'd5839: data = 8'h1b;
      17'd5840: data = 8'h22;
      17'd5841: data = 8'h19;
      17'd5842: data = 8'h16;
      17'd5843: data = 8'h1b;
      17'd5844: data = 8'h1b;
      17'd5845: data = 8'h16;
      17'd5846: data = 8'h11;
      17'd5847: data = 8'h16;
      17'd5848: data = 8'h13;
      17'd5849: data = 8'h11;
      17'd5850: data = 8'h13;
      17'd5851: data = 8'h09;
      17'd5852: data = 8'h0a;
      17'd5853: data = 8'h0d;
      17'd5854: data = 8'h02;
      17'd5855: data = 8'hfd;
      17'd5856: data = 8'h00;
      17'd5857: data = 8'h06;
      17'd5858: data = 8'hfe;
      17'd5859: data = 8'hf5;
      17'd5860: data = 8'hf9;
      17'd5861: data = 8'hf9;
      17'd5862: data = 8'hf6;
      17'd5863: data = 8'hfa;
      17'd5864: data = 8'hf9;
      17'd5865: data = 8'hf1;
      17'd5866: data = 8'hed;
      17'd5867: data = 8'hf1;
      17'd5868: data = 8'hf2;
      17'd5869: data = 8'hf2;
      17'd5870: data = 8'hf2;
      17'd5871: data = 8'hef;
      17'd5872: data = 8'hef;
      17'd5873: data = 8'hf2;
      17'd5874: data = 8'hf4;
      17'd5875: data = 8'hf4;
      17'd5876: data = 8'hf4;
      17'd5877: data = 8'hfc;
      17'd5878: data = 8'hfc;
      17'd5879: data = 8'hfd;
      17'd5880: data = 8'hfd;
      17'd5881: data = 8'hfc;
      17'd5882: data = 8'h01;
      17'd5883: data = 8'h02;
      17'd5884: data = 8'h01;
      17'd5885: data = 8'h09;
      17'd5886: data = 8'h0c;
      17'd5887: data = 8'h0d;
      17'd5888: data = 8'h0d;
      17'd5889: data = 8'h0e;
      17'd5890: data = 8'h11;
      17'd5891: data = 8'h0e;
      17'd5892: data = 8'h15;
      17'd5893: data = 8'h1b;
      17'd5894: data = 8'h1a;
      17'd5895: data = 8'h1c;
      17'd5896: data = 8'h1c;
      17'd5897: data = 8'h1a;
      17'd5898: data = 8'h1b;
      17'd5899: data = 8'h19;
      17'd5900: data = 8'h0e;
      17'd5901: data = 8'h16;
      17'd5902: data = 8'h1f;
      17'd5903: data = 8'h22;
      17'd5904: data = 8'h26;
      17'd5905: data = 8'h26;
      17'd5906: data = 8'h22;
      17'd5907: data = 8'h1e;
      17'd5908: data = 8'h15;
      17'd5909: data = 8'h15;
      17'd5910: data = 8'h1b;
      17'd5911: data = 8'h16;
      17'd5912: data = 8'h16;
      17'd5913: data = 8'h1c;
      17'd5914: data = 8'h1a;
      17'd5915: data = 8'h1c;
      17'd5916: data = 8'h15;
      17'd5917: data = 8'h0d;
      17'd5918: data = 8'h11;
      17'd5919: data = 8'h13;
      17'd5920: data = 8'h12;
      17'd5921: data = 8'h0a;
      17'd5922: data = 8'h09;
      17'd5923: data = 8'h12;
      17'd5924: data = 8'h0d;
      17'd5925: data = 8'h00;
      17'd5926: data = 8'hfe;
      17'd5927: data = 8'h04;
      17'd5928: data = 8'h04;
      17'd5929: data = 8'hfa;
      17'd5930: data = 8'hfe;
      17'd5931: data = 8'h00;
      17'd5932: data = 8'hf4;
      17'd5933: data = 8'hef;
      17'd5934: data = 8'hf1;
      17'd5935: data = 8'hec;
      17'd5936: data = 8'he7;
      17'd5937: data = 8'hed;
      17'd5938: data = 8'he9;
      17'd5939: data = 8'he4;
      17'd5940: data = 8'he5;
      17'd5941: data = 8'he2;
      17'd5942: data = 8'hd8;
      17'd5943: data = 8'hd6;
      17'd5944: data = 8'hd5;
      17'd5945: data = 8'hd3;
      17'd5946: data = 8'hd1;
      17'd5947: data = 8'hd2;
      17'd5948: data = 8'hd2;
      17'd5949: data = 8'hcb;
      17'd5950: data = 8'hcd;
      17'd5951: data = 8'hcd;
      17'd5952: data = 8'hc5;
      17'd5953: data = 8'hc4;
      17'd5954: data = 8'hc6;
      17'd5955: data = 8'hc4;
      17'd5956: data = 8'hc9;
      17'd5957: data = 8'hc9;
      17'd5958: data = 8'hc4;
      17'd5959: data = 8'hc4;
      17'd5960: data = 8'hc6;
      17'd5961: data = 8'hc6;
      17'd5962: data = 8'hc6;
      17'd5963: data = 8'hc9;
      17'd5964: data = 8'hd1;
      17'd5965: data = 8'hd5;
      17'd5966: data = 8'hcb;
      17'd5967: data = 8'hc9;
      17'd5968: data = 8'hd2;
      17'd5969: data = 8'he2;
      17'd5970: data = 8'hdb;
      17'd5971: data = 8'hdb;
      17'd5972: data = 8'he7;
      17'd5973: data = 8'he5;
      17'd5974: data = 8'he7;
      17'd5975: data = 8'hf1;
      17'd5976: data = 8'hf5;
      17'd5977: data = 8'hed;
      17'd5978: data = 8'hec;
      17'd5979: data = 8'hf5;
      17'd5980: data = 8'h01;
      17'd5981: data = 8'hfe;
      17'd5982: data = 8'h04;
      17'd5983: data = 8'h06;
      17'd5984: data = 8'hfe;
      17'd5985: data = 8'h02;
      17'd5986: data = 8'h15;
      17'd5987: data = 8'h12;
      17'd5988: data = 8'h09;
      17'd5989: data = 8'h11;
      17'd5990: data = 8'h16;
      17'd5991: data = 8'h0e;
      17'd5992: data = 8'hfd;
      17'd5993: data = 8'h1f;
      17'd5994: data = 8'h1a;
      17'd5995: data = 8'h0a;
      17'd5996: data = 8'h22;
      17'd5997: data = 8'h15;
      17'd5998: data = 8'h13;
      17'd5999: data = 8'h11;
      17'd6000: data = 8'h16;
      17'd6001: data = 8'h1a;
      17'd6002: data = 8'h06;
      17'd6003: data = 8'h12;
      17'd6004: data = 8'h12;
      17'd6005: data = 8'h0c;
      17'd6006: data = 8'h1a;
      17'd6007: data = 8'h16;
      17'd6008: data = 8'h13;
      17'd6009: data = 8'h05;
      17'd6010: data = 8'h01;
      17'd6011: data = 8'hfe;
      17'd6012: data = 8'hf6;
      17'd6013: data = 8'hfe;
      17'd6014: data = 8'h04;
      17'd6015: data = 8'h0a;
      17'd6016: data = 8'h0a;
      17'd6017: data = 8'hfe;
      17'd6018: data = 8'hf9;
      17'd6019: data = 8'hfe;
      17'd6020: data = 8'hfa;
      17'd6021: data = 8'hf6;
      17'd6022: data = 8'h0d;
      17'd6023: data = 8'h09;
      17'd6024: data = 8'hf5;
      17'd6025: data = 8'hfd;
      17'd6026: data = 8'h00;
      17'd6027: data = 8'hf2;
      17'd6028: data = 8'hf9;
      17'd6029: data = 8'h06;
      17'd6030: data = 8'h0a;
      17'd6031: data = 8'h0e;
      17'd6032: data = 8'h0d;
      17'd6033: data = 8'h06;
      17'd6034: data = 8'h05;
      17'd6035: data = 8'h05;
      17'd6036: data = 8'h09;
      17'd6037: data = 8'h05;
      17'd6038: data = 8'h06;
      17'd6039: data = 8'h12;
      17'd6040: data = 8'h19;
      17'd6041: data = 8'h12;
      17'd6042: data = 8'h0e;
      17'd6043: data = 8'h1a;
      17'd6044: data = 8'h1e;
      17'd6045: data = 8'h13;
      17'd6046: data = 8'h15;
      17'd6047: data = 8'h1c;
      17'd6048: data = 8'h15;
      17'd6049: data = 8'h11;
      17'd6050: data = 8'h1a;
      17'd6051: data = 8'h1e;
      17'd6052: data = 8'h1b;
      17'd6053: data = 8'h1b;
      17'd6054: data = 8'h1b;
      17'd6055: data = 8'h16;
      17'd6056: data = 8'h16;
      17'd6057: data = 8'h1c;
      17'd6058: data = 8'h1c;
      17'd6059: data = 8'h1a;
      17'd6060: data = 8'h16;
      17'd6061: data = 8'h13;
      17'd6062: data = 8'h0d;
      17'd6063: data = 8'h04;
      17'd6064: data = 8'h0d;
      17'd6065: data = 8'h12;
      17'd6066: data = 8'h06;
      17'd6067: data = 8'h0e;
      17'd6068: data = 8'h13;
      17'd6069: data = 8'h01;
      17'd6070: data = 8'hfd;
      17'd6071: data = 8'h01;
      17'd6072: data = 8'hfd;
      17'd6073: data = 8'hf9;
      17'd6074: data = 8'hfc;
      17'd6075: data = 8'hfd;
      17'd6076: data = 8'hfc;
      17'd6077: data = 8'hfa;
      17'd6078: data = 8'hfa;
      17'd6079: data = 8'hfa;
      17'd6080: data = 8'hf5;
      17'd6081: data = 8'hf5;
      17'd6082: data = 8'hf4;
      17'd6083: data = 8'hf2;
      17'd6084: data = 8'hf1;
      17'd6085: data = 8'hf6;
      17'd6086: data = 8'hf6;
      17'd6087: data = 8'hf4;
      17'd6088: data = 8'hf6;
      17'd6089: data = 8'hf9;
      17'd6090: data = 8'hfa;
      17'd6091: data = 8'hfa;
      17'd6092: data = 8'hfa;
      17'd6093: data = 8'hfc;
      17'd6094: data = 8'hfd;
      17'd6095: data = 8'hfe;
      17'd6096: data = 8'h00;
      17'd6097: data = 8'h01;
      17'd6098: data = 8'h00;
      17'd6099: data = 8'h01;
      17'd6100: data = 8'h04;
      17'd6101: data = 8'h05;
      17'd6102: data = 8'h09;
      17'd6103: data = 8'h11;
      17'd6104: data = 8'h12;
      17'd6105: data = 8'h0d;
      17'd6106: data = 8'h0e;
      17'd6107: data = 8'h0c;
      17'd6108: data = 8'h0d;
      17'd6109: data = 8'h11;
      17'd6110: data = 8'h11;
      17'd6111: data = 8'h13;
      17'd6112: data = 8'h15;
      17'd6113: data = 8'h13;
      17'd6114: data = 8'h15;
      17'd6115: data = 8'h13;
      17'd6116: data = 8'h15;
      17'd6117: data = 8'h15;
      17'd6118: data = 8'h15;
      17'd6119: data = 8'h1a;
      17'd6120: data = 8'h16;
      17'd6121: data = 8'h13;
      17'd6122: data = 8'h0e;
      17'd6123: data = 8'h12;
      17'd6124: data = 8'h1a;
      17'd6125: data = 8'h13;
      17'd6126: data = 8'h0d;
      17'd6127: data = 8'h15;
      17'd6128: data = 8'h19;
      17'd6129: data = 8'h11;
      17'd6130: data = 8'h0e;
      17'd6131: data = 8'h0d;
      17'd6132: data = 8'h0c;
      17'd6133: data = 8'h0a;
      17'd6134: data = 8'h09;
      17'd6135: data = 8'h0c;
      17'd6136: data = 8'h09;
      17'd6137: data = 8'h06;
      17'd6138: data = 8'h0a;
      17'd6139: data = 8'h04;
      17'd6140: data = 8'h01;
      17'd6141: data = 8'h01;
      17'd6142: data = 8'hfd;
      17'd6143: data = 8'hfd;
      17'd6144: data = 8'hfc;
      17'd6145: data = 8'hf6;
      17'd6146: data = 8'hf5;
      17'd6147: data = 8'hf2;
      17'd6148: data = 8'hf1;
      17'd6149: data = 8'hed;
      17'd6150: data = 8'hed;
      17'd6151: data = 8'heb;
      17'd6152: data = 8'he4;
      17'd6153: data = 8'he5;
      17'd6154: data = 8'he2;
      17'd6155: data = 8'he0;
      17'd6156: data = 8'hde;
      17'd6157: data = 8'hdb;
      17'd6158: data = 8'hd8;
      17'd6159: data = 8'hd3;
      17'd6160: data = 8'hd6;
      17'd6161: data = 8'hd3;
      17'd6162: data = 8'hd2;
      17'd6163: data = 8'hd6;
      17'd6164: data = 8'hcd;
      17'd6165: data = 8'hc6;
      17'd6166: data = 8'hce;
      17'd6167: data = 8'hd2;
      17'd6168: data = 8'hc6;
      17'd6169: data = 8'hc6;
      17'd6170: data = 8'hcb;
      17'd6171: data = 8'hca;
      17'd6172: data = 8'hcb;
      17'd6173: data = 8'hd1;
      17'd6174: data = 8'hd1;
      17'd6175: data = 8'hce;
      17'd6176: data = 8'hcb;
      17'd6177: data = 8'hcd;
      17'd6178: data = 8'hd3;
      17'd6179: data = 8'hd3;
      17'd6180: data = 8'hda;
      17'd6181: data = 8'hdc;
      17'd6182: data = 8'hde;
      17'd6183: data = 8'he3;
      17'd6184: data = 8'he0;
      17'd6185: data = 8'hdc;
      17'd6186: data = 8'hec;
      17'd6187: data = 8'hf1;
      17'd6188: data = 8'heb;
      17'd6189: data = 8'hec;
      17'd6190: data = 8'hf4;
      17'd6191: data = 8'hfd;
      17'd6192: data = 8'hf4;
      17'd6193: data = 8'hf9;
      17'd6194: data = 8'h04;
      17'd6195: data = 8'h01;
      17'd6196: data = 8'h04;
      17'd6197: data = 8'h04;
      17'd6198: data = 8'h0a;
      17'd6199: data = 8'h05;
      17'd6200: data = 8'h09;
      17'd6201: data = 8'h0e;
      17'd6202: data = 8'h0a;
      17'd6203: data = 8'h0e;
      17'd6204: data = 8'h1c;
      17'd6205: data = 8'h12;
      17'd6206: data = 8'h0e;
      17'd6207: data = 8'h19;
      17'd6208: data = 8'h19;
      17'd6209: data = 8'h12;
      17'd6210: data = 8'h15;
      17'd6211: data = 8'h1a;
      17'd6212: data = 8'h0a;
      17'd6213: data = 8'h13;
      17'd6214: data = 8'h1c;
      17'd6215: data = 8'h16;
      17'd6216: data = 8'h16;
      17'd6217: data = 8'h0e;
      17'd6218: data = 8'h0c;
      17'd6219: data = 8'h0e;
      17'd6220: data = 8'h11;
      17'd6221: data = 8'h12;
      17'd6222: data = 8'h0e;
      17'd6223: data = 8'h0a;
      17'd6224: data = 8'hfe;
      17'd6225: data = 8'hfa;
      17'd6226: data = 8'hfd;
      17'd6227: data = 8'hf6;
      17'd6228: data = 8'h00;
      17'd6229: data = 8'h06;
      17'd6230: data = 8'h00;
      17'd6231: data = 8'h04;
      17'd6232: data = 8'h01;
      17'd6233: data = 8'hf4;
      17'd6234: data = 8'hfd;
      17'd6235: data = 8'h04;
      17'd6236: data = 8'h01;
      17'd6237: data = 8'hfe;
      17'd6238: data = 8'h00;
      17'd6239: data = 8'hfa;
      17'd6240: data = 8'hef;
      17'd6241: data = 8'hfc;
      17'd6242: data = 8'h02;
      17'd6243: data = 8'h05;
      17'd6244: data = 8'h0d;
      17'd6245: data = 8'h0e;
      17'd6246: data = 8'h09;
      17'd6247: data = 8'h00;
      17'd6248: data = 8'h02;
      17'd6249: data = 8'h06;
      17'd6250: data = 8'h0c;
      17'd6251: data = 8'h12;
      17'd6252: data = 8'h12;
      17'd6253: data = 8'h12;
      17'd6254: data = 8'h13;
      17'd6255: data = 8'h0d;
      17'd6256: data = 8'h15;
      17'd6257: data = 8'h1c;
      17'd6258: data = 8'h19;
      17'd6259: data = 8'h1a;
      17'd6260: data = 8'h1a;
      17'd6261: data = 8'h15;
      17'd6262: data = 8'h13;
      17'd6263: data = 8'h15;
      17'd6264: data = 8'h1b;
      17'd6265: data = 8'h1e;
      17'd6266: data = 8'h22;
      17'd6267: data = 8'h23;
      17'd6268: data = 8'h1b;
      17'd6269: data = 8'h1a;
      17'd6270: data = 8'h19;
      17'd6271: data = 8'h16;
      17'd6272: data = 8'h13;
      17'd6273: data = 8'h12;
      17'd6274: data = 8'h13;
      17'd6275: data = 8'h11;
      17'd6276: data = 8'h0c;
      17'd6277: data = 8'h0c;
      17'd6278: data = 8'h0d;
      17'd6279: data = 8'h09;
      17'd6280: data = 8'h06;
      17'd6281: data = 8'h0c;
      17'd6282: data = 8'h06;
      17'd6283: data = 8'h00;
      17'd6284: data = 8'h00;
      17'd6285: data = 8'hfd;
      17'd6286: data = 8'hfc;
      17'd6287: data = 8'hf9;
      17'd6288: data = 8'hf9;
      17'd6289: data = 8'hfc;
      17'd6290: data = 8'hf5;
      17'd6291: data = 8'hf9;
      17'd6292: data = 8'hf9;
      17'd6293: data = 8'hf6;
      17'd6294: data = 8'hf6;
      17'd6295: data = 8'hf5;
      17'd6296: data = 8'hf5;
      17'd6297: data = 8'hf6;
      17'd6298: data = 8'hf2;
      17'd6299: data = 8'hf2;
      17'd6300: data = 8'hf2;
      17'd6301: data = 8'hf5;
      17'd6302: data = 8'hfd;
      17'd6303: data = 8'hfc;
      17'd6304: data = 8'hfd;
      17'd6305: data = 8'hfc;
      17'd6306: data = 8'hfc;
      17'd6307: data = 8'hfa;
      17'd6308: data = 8'hfc;
      17'd6309: data = 8'h01;
      17'd6310: data = 8'h02;
      17'd6311: data = 8'h01;
      17'd6312: data = 8'hfe;
      17'd6313: data = 8'h02;
      17'd6314: data = 8'h09;
      17'd6315: data = 8'h09;
      17'd6316: data = 8'h0a;
      17'd6317: data = 8'h11;
      17'd6318: data = 8'h0d;
      17'd6319: data = 8'h0c;
      17'd6320: data = 8'h0d;
      17'd6321: data = 8'h0c;
      17'd6322: data = 8'h0e;
      17'd6323: data = 8'h0e;
      17'd6324: data = 8'h0a;
      17'd6325: data = 8'h11;
      17'd6326: data = 8'h15;
      17'd6327: data = 8'h11;
      17'd6328: data = 8'h11;
      17'd6329: data = 8'h12;
      17'd6330: data = 8'h12;
      17'd6331: data = 8'h0c;
      17'd6332: data = 8'h0c;
      17'd6333: data = 8'h12;
      17'd6334: data = 8'h0d;
      17'd6335: data = 8'h0e;
      17'd6336: data = 8'h13;
      17'd6337: data = 8'h0d;
      17'd6338: data = 8'h0c;
      17'd6339: data = 8'h11;
      17'd6340: data = 8'h0d;
      17'd6341: data = 8'h09;
      17'd6342: data = 8'h0a;
      17'd6343: data = 8'h09;
      17'd6344: data = 8'h06;
      17'd6345: data = 8'h04;
      17'd6346: data = 8'h04;
      17'd6347: data = 8'h05;
      17'd6348: data = 8'h01;
      17'd6349: data = 8'hfe;
      17'd6350: data = 8'h01;
      17'd6351: data = 8'h02;
      17'd6352: data = 8'hfe;
      17'd6353: data = 8'hfd;
      17'd6354: data = 8'hfe;
      17'd6355: data = 8'hfd;
      17'd6356: data = 8'hfa;
      17'd6357: data = 8'hfa;
      17'd6358: data = 8'hf6;
      17'd6359: data = 8'hfa;
      17'd6360: data = 8'hf9;
      17'd6361: data = 8'hef;
      17'd6362: data = 8'hef;
      17'd6363: data = 8'hf6;
      17'd6364: data = 8'hf2;
      17'd6365: data = 8'hec;
      17'd6366: data = 8'hf2;
      17'd6367: data = 8'hf1;
      17'd6368: data = 8'hec;
      17'd6369: data = 8'heb;
      17'd6370: data = 8'heb;
      17'd6371: data = 8'hec;
      17'd6372: data = 8'he9;
      17'd6373: data = 8'he5;
      17'd6374: data = 8'he7;
      17'd6375: data = 8'heb;
      17'd6376: data = 8'he7;
      17'd6377: data = 8'he3;
      17'd6378: data = 8'he3;
      17'd6379: data = 8'he2;
      17'd6380: data = 8'he3;
      17'd6381: data = 8'he2;
      17'd6382: data = 8'hde;
      17'd6383: data = 8'hdc;
      17'd6384: data = 8'hda;
      17'd6385: data = 8'hdb;
      17'd6386: data = 8'hdb;
      17'd6387: data = 8'he0;
      17'd6388: data = 8'he0;
      17'd6389: data = 8'hdb;
      17'd6390: data = 8'hde;
      17'd6391: data = 8'hde;
      17'd6392: data = 8'hdb;
      17'd6393: data = 8'hdc;
      17'd6394: data = 8'hdc;
      17'd6395: data = 8'hdc;
      17'd6396: data = 8'he2;
      17'd6397: data = 8'hde;
      17'd6398: data = 8'hdc;
      17'd6399: data = 8'he2;
      17'd6400: data = 8'he2;
      17'd6401: data = 8'he5;
      17'd6402: data = 8'he9;
      17'd6403: data = 8'he5;
      17'd6404: data = 8'heb;
      17'd6405: data = 8'hed;
      17'd6406: data = 8'heb;
      17'd6407: data = 8'hed;
      17'd6408: data = 8'hef;
      17'd6409: data = 8'hf2;
      17'd6410: data = 8'hf5;
      17'd6411: data = 8'hf6;
      17'd6412: data = 8'hf9;
      17'd6413: data = 8'hfa;
      17'd6414: data = 8'hfc;
      17'd6415: data = 8'h00;
      17'd6416: data = 8'h04;
      17'd6417: data = 8'h04;
      17'd6418: data = 8'h09;
      17'd6419: data = 8'h0c;
      17'd6420: data = 8'h09;
      17'd6421: data = 8'h06;
      17'd6422: data = 8'h0d;
      17'd6423: data = 8'h11;
      17'd6424: data = 8'h0e;
      17'd6425: data = 8'h0e;
      17'd6426: data = 8'h11;
      17'd6427: data = 8'h12;
      17'd6428: data = 8'h13;
      17'd6429: data = 8'h16;
      17'd6430: data = 8'h15;
      17'd6431: data = 8'h16;
      17'd6432: data = 8'h1b;
      17'd6433: data = 8'h19;
      17'd6434: data = 8'h15;
      17'd6435: data = 8'h16;
      17'd6436: data = 8'h15;
      17'd6437: data = 8'h13;
      17'd6438: data = 8'h15;
      17'd6439: data = 8'h16;
      17'd6440: data = 8'h15;
      17'd6441: data = 8'h13;
      17'd6442: data = 8'h19;
      17'd6443: data = 8'h19;
      17'd6444: data = 8'h15;
      17'd6445: data = 8'h13;
      17'd6446: data = 8'h12;
      17'd6447: data = 8'h12;
      17'd6448: data = 8'h15;
      17'd6449: data = 8'h12;
      17'd6450: data = 8'h0e;
      17'd6451: data = 8'h0c;
      17'd6452: data = 8'h0d;
      17'd6453: data = 8'h0d;
      17'd6454: data = 8'h0c;
      17'd6455: data = 8'h0a;
      17'd6456: data = 8'h0c;
      17'd6457: data = 8'h0c;
      17'd6458: data = 8'h06;
      17'd6459: data = 8'h04;
      17'd6460: data = 8'h09;
      17'd6461: data = 8'h0a;
      17'd6462: data = 8'h09;
      17'd6463: data = 8'h06;
      17'd6464: data = 8'h01;
      17'd6465: data = 8'h04;
      17'd6466: data = 8'h06;
      17'd6467: data = 8'h04;
      17'd6468: data = 8'h04;
      17'd6469: data = 8'h02;
      17'd6470: data = 8'h01;
      17'd6471: data = 8'h01;
      17'd6472: data = 8'h04;
      17'd6473: data = 8'h02;
      17'd6474: data = 8'h00;
      17'd6475: data = 8'h00;
      17'd6476: data = 8'h05;
      17'd6477: data = 8'h09;
      17'd6478: data = 8'h02;
      17'd6479: data = 8'hfe;
      17'd6480: data = 8'h06;
      17'd6481: data = 8'h0c;
      17'd6482: data = 8'h06;
      17'd6483: data = 8'h04;
      17'd6484: data = 8'h05;
      17'd6485: data = 8'h0a;
      17'd6486: data = 8'h0a;
      17'd6487: data = 8'h09;
      17'd6488: data = 8'h09;
      17'd6489: data = 8'h09;
      17'd6490: data = 8'h0d;
      17'd6491: data = 8'h0e;
      17'd6492: data = 8'h0a;
      17'd6493: data = 8'h06;
      17'd6494: data = 8'h0a;
      17'd6495: data = 8'h09;
      17'd6496: data = 8'h0a;
      17'd6497: data = 8'h09;
      17'd6498: data = 8'h06;
      17'd6499: data = 8'h06;
      17'd6500: data = 8'h09;
      17'd6501: data = 8'h06;
      17'd6502: data = 8'h06;
      17'd6503: data = 8'h05;
      17'd6504: data = 8'h00;
      17'd6505: data = 8'h02;
      17'd6506: data = 8'h05;
      17'd6507: data = 8'h02;
      17'd6508: data = 8'hfd;
      17'd6509: data = 8'hfe;
      17'd6510: data = 8'h01;
      17'd6511: data = 8'h00;
      17'd6512: data = 8'h01;
      17'd6513: data = 8'hfa;
      17'd6514: data = 8'hf9;
      17'd6515: data = 8'hfd;
      17'd6516: data = 8'hfa;
      17'd6517: data = 8'hfa;
      17'd6518: data = 8'hfa;
      17'd6519: data = 8'hf9;
      17'd6520: data = 8'hf5;
      17'd6521: data = 8'hf4;
      17'd6522: data = 8'hf4;
      17'd6523: data = 8'hf4;
      17'd6524: data = 8'hf5;
      17'd6525: data = 8'hf6;
      17'd6526: data = 8'hfa;
      17'd6527: data = 8'hf5;
      17'd6528: data = 8'hf5;
      17'd6529: data = 8'hf9;
      17'd6530: data = 8'hf6;
      17'd6531: data = 8'hf5;
      17'd6532: data = 8'hf5;
      17'd6533: data = 8'hfc;
      17'd6534: data = 8'hf4;
      17'd6535: data = 8'hf2;
      17'd6536: data = 8'hf9;
      17'd6537: data = 8'hf6;
      17'd6538: data = 8'hf5;
      17'd6539: data = 8'hf5;
      17'd6540: data = 8'hf9;
      17'd6541: data = 8'hf9;
      17'd6542: data = 8'hfa;
      17'd6543: data = 8'hfc;
      17'd6544: data = 8'hfa;
      17'd6545: data = 8'hf6;
      17'd6546: data = 8'hf9;
      17'd6547: data = 8'hfa;
      17'd6548: data = 8'hfc;
      17'd6549: data = 8'hfa;
      17'd6550: data = 8'hf6;
      17'd6551: data = 8'hfa;
      17'd6552: data = 8'hfc;
      17'd6553: data = 8'hf9;
      17'd6554: data = 8'hfc;
      17'd6555: data = 8'hf9;
      17'd6556: data = 8'hf9;
      17'd6557: data = 8'hfd;
      17'd6558: data = 8'hf6;
      17'd6559: data = 8'hf9;
      17'd6560: data = 8'hfe;
      17'd6561: data = 8'hfc;
      17'd6562: data = 8'hf9;
      17'd6563: data = 8'hfc;
      17'd6564: data = 8'hfe;
      17'd6565: data = 8'hfc;
      17'd6566: data = 8'hfd;
      17'd6567: data = 8'hfe;
      17'd6568: data = 8'hfd;
      17'd6569: data = 8'hfc;
      17'd6570: data = 8'hfc;
      17'd6571: data = 8'hfd;
      17'd6572: data = 8'hfd;
      17'd6573: data = 8'h00;
      17'd6574: data = 8'h00;
      17'd6575: data = 8'hfc;
      17'd6576: data = 8'hfd;
      17'd6577: data = 8'h01;
      17'd6578: data = 8'h01;
      17'd6579: data = 8'hfd;
      17'd6580: data = 8'hfd;
      17'd6581: data = 8'h01;
      17'd6582: data = 8'hfd;
      17'd6583: data = 8'hfd;
      17'd6584: data = 8'hfe;
      17'd6585: data = 8'hfd;
      17'd6586: data = 8'hfe;
      17'd6587: data = 8'hfc;
      17'd6588: data = 8'hf9;
      17'd6589: data = 8'hfc;
      17'd6590: data = 8'hfa;
      17'd6591: data = 8'hfa;
      17'd6592: data = 8'hfa;
      17'd6593: data = 8'hf6;
      17'd6594: data = 8'hfa;
      17'd6595: data = 8'hfa;
      17'd6596: data = 8'hf9;
      17'd6597: data = 8'hfc;
      17'd6598: data = 8'hf9;
      17'd6599: data = 8'hf4;
      17'd6600: data = 8'hf6;
      17'd6601: data = 8'hf9;
      17'd6602: data = 8'hf6;
      17'd6603: data = 8'hf4;
      17'd6604: data = 8'hf4;
      17'd6605: data = 8'hf6;
      17'd6606: data = 8'hf5;
      17'd6607: data = 8'hf4;
      17'd6608: data = 8'hf5;
      17'd6609: data = 8'hf6;
      17'd6610: data = 8'hf2;
      17'd6611: data = 8'hf5;
      17'd6612: data = 8'hf6;
      17'd6613: data = 8'hf4;
      17'd6614: data = 8'hf4;
      17'd6615: data = 8'hf6;
      17'd6616: data = 8'hf5;
      17'd6617: data = 8'hf6;
      17'd6618: data = 8'hf4;
      17'd6619: data = 8'hf1;
      17'd6620: data = 8'hf4;
      17'd6621: data = 8'hf6;
      17'd6622: data = 8'hf6;
      17'd6623: data = 8'hf4;
      17'd6624: data = 8'hf4;
      17'd6625: data = 8'hfc;
      17'd6626: data = 8'hf9;
      17'd6627: data = 8'hfa;
      17'd6628: data = 8'hfc;
      17'd6629: data = 8'hf9;
      17'd6630: data = 8'hfc;
      17'd6631: data = 8'hfa;
      17'd6632: data = 8'hf9;
      17'd6633: data = 8'hfc;
      17'd6634: data = 8'hfc;
      17'd6635: data = 8'hfd;
      17'd6636: data = 8'hfc;
      17'd6637: data = 8'hf9;
      17'd6638: data = 8'hfc;
      17'd6639: data = 8'h00;
      17'd6640: data = 8'h00;
      17'd6641: data = 8'h00;
      17'd6642: data = 8'hfd;
      17'd6643: data = 8'hfe;
      17'd6644: data = 8'hfe;
      17'd6645: data = 8'h01;
      17'd6646: data = 8'h01;
      17'd6647: data = 8'hfc;
      17'd6648: data = 8'hfe;
      17'd6649: data = 8'h02;
      17'd6650: data = 8'hfe;
      17'd6651: data = 8'h00;
      17'd6652: data = 8'h01;
      17'd6653: data = 8'h02;
      17'd6654: data = 8'h02;
      17'd6655: data = 8'h05;
      17'd6656: data = 8'h02;
      17'd6657: data = 8'h01;
      17'd6658: data = 8'h09;
      17'd6659: data = 8'h05;
      17'd6660: data = 8'h04;
      17'd6661: data = 8'h05;
      17'd6662: data = 8'h05;
      17'd6663: data = 8'h09;
      17'd6664: data = 8'h09;
      17'd6665: data = 8'h0c;
      17'd6666: data = 8'h0c;
      17'd6667: data = 8'h05;
      17'd6668: data = 8'h09;
      17'd6669: data = 8'h0d;
      17'd6670: data = 8'h0c;
      17'd6671: data = 8'h0c;
      17'd6672: data = 8'h0c;
      17'd6673: data = 8'h0c;
      17'd6674: data = 8'h0e;
      17'd6675: data = 8'h0e;
      17'd6676: data = 8'h0d;
      17'd6677: data = 8'h0e;
      17'd6678: data = 8'h0e;
      17'd6679: data = 8'h0d;
      17'd6680: data = 8'h0d;
      17'd6681: data = 8'h0e;
      17'd6682: data = 8'h0d;
      17'd6683: data = 8'h0e;
      17'd6684: data = 8'h0d;
      17'd6685: data = 8'h0c;
      17'd6686: data = 8'h0c;
      17'd6687: data = 8'h0c;
      17'd6688: data = 8'h0c;
      17'd6689: data = 8'h0c;
      17'd6690: data = 8'h0c;
      17'd6691: data = 8'h0c;
      17'd6692: data = 8'h09;
      17'd6693: data = 8'h06;
      17'd6694: data = 8'h0c;
      17'd6695: data = 8'h0a;
      17'd6696: data = 8'h04;
      17'd6697: data = 8'h05;
      17'd6698: data = 8'h0a;
      17'd6699: data = 8'h06;
      17'd6700: data = 8'h06;
      17'd6701: data = 8'h06;
      17'd6702: data = 8'h0a;
      17'd6703: data = 8'h09;
      17'd6704: data = 8'h04;
      17'd6705: data = 8'h02;
      17'd6706: data = 8'h04;
      17'd6707: data = 8'h02;
      17'd6708: data = 8'h00;
      17'd6709: data = 8'h00;
      17'd6710: data = 8'h00;
      17'd6711: data = 8'h00;
      17'd6712: data = 8'h00;
      17'd6713: data = 8'hfc;
      17'd6714: data = 8'hfe;
      17'd6715: data = 8'h00;
      17'd6716: data = 8'hfc;
      17'd6717: data = 8'hfd;
      17'd6718: data = 8'hfc;
      17'd6719: data = 8'hfc;
      17'd6720: data = 8'hfc;
      17'd6721: data = 8'hfa;
      17'd6722: data = 8'hfa;
      17'd6723: data = 8'hfa;
      17'd6724: data = 8'hfc;
      17'd6725: data = 8'hf9;
      17'd6726: data = 8'hfc;
      17'd6727: data = 8'hfd;
      17'd6728: data = 8'hfa;
      17'd6729: data = 8'hf9;
      17'd6730: data = 8'hf9;
      17'd6731: data = 8'hfa;
      17'd6732: data = 8'hfc;
      17'd6733: data = 8'hfa;
      17'd6734: data = 8'hf9;
      17'd6735: data = 8'hfa;
      17'd6736: data = 8'hfa;
      17'd6737: data = 8'hf9;
      17'd6738: data = 8'hfc;
      17'd6739: data = 8'hfc;
      17'd6740: data = 8'hfc;
      17'd6741: data = 8'hfc;
      17'd6742: data = 8'hfd;
      17'd6743: data = 8'hfd;
      17'd6744: data = 8'hfc;
      17'd6745: data = 8'hfe;
      17'd6746: data = 8'hfc;
      17'd6747: data = 8'hfc;
      17'd6748: data = 8'hfc;
      17'd6749: data = 8'hfc;
      17'd6750: data = 8'hfe;
      17'd6751: data = 8'hfe;
      17'd6752: data = 8'hfc;
      17'd6753: data = 8'hfc;
      17'd6754: data = 8'hfc;
      17'd6755: data = 8'hfc;
      17'd6756: data = 8'h00;
      17'd6757: data = 8'hfd;
      17'd6758: data = 8'hfa;
      17'd6759: data = 8'hfd;
      17'd6760: data = 8'hf9;
      17'd6761: data = 8'hfc;
      17'd6762: data = 8'hfc;
      17'd6763: data = 8'hf6;
      17'd6764: data = 8'hfe;
      17'd6765: data = 8'h00;
      17'd6766: data = 8'hf9;
      17'd6767: data = 8'hfd;
      17'd6768: data = 8'hfe;
      17'd6769: data = 8'hfa;
      17'd6770: data = 8'hfc;
      17'd6771: data = 8'hfd;
      17'd6772: data = 8'hfa;
      17'd6773: data = 8'hfc;
      17'd6774: data = 8'hfd;
      17'd6775: data = 8'hfc;
      17'd6776: data = 8'hf9;
      17'd6777: data = 8'hfe;
      17'd6778: data = 8'h01;
      17'd6779: data = 8'hfe;
      17'd6780: data = 8'hfd;
      17'd6781: data = 8'h01;
      17'd6782: data = 8'h04;
      17'd6783: data = 8'h00;
      17'd6784: data = 8'hfc;
      17'd6785: data = 8'hfe;
      17'd6786: data = 8'h02;
      17'd6787: data = 8'hfe;
      17'd6788: data = 8'hfd;
      17'd6789: data = 8'h00;
      17'd6790: data = 8'h01;
      17'd6791: data = 8'h02;
      17'd6792: data = 8'h02;
      17'd6793: data = 8'h02;
      17'd6794: data = 8'h06;
      17'd6795: data = 8'h04;
      17'd6796: data = 8'h02;
      17'd6797: data = 8'h04;
      17'd6798: data = 8'h01;
      17'd6799: data = 8'h01;
      17'd6800: data = 8'h00;
      17'd6801: data = 8'h02;
      17'd6802: data = 8'h04;
      17'd6803: data = 8'h04;
      17'd6804: data = 8'h04;
      17'd6805: data = 8'h02;
      17'd6806: data = 8'h04;
      17'd6807: data = 8'h05;
      17'd6808: data = 8'h04;
      17'd6809: data = 8'h01;
      17'd6810: data = 8'h01;
      17'd6811: data = 8'h02;
      17'd6812: data = 8'h02;
      17'd6813: data = 8'h00;
      17'd6814: data = 8'h01;
      17'd6815: data = 8'h01;
      17'd6816: data = 8'hfd;
      17'd6817: data = 8'h00;
      17'd6818: data = 8'h02;
      17'd6819: data = 8'h00;
      17'd6820: data = 8'hfd;
      17'd6821: data = 8'hfe;
      17'd6822: data = 8'h01;
      17'd6823: data = 8'h01;
      17'd6824: data = 8'hfd;
      17'd6825: data = 8'h00;
      17'd6826: data = 8'h00;
      17'd6827: data = 8'hfd;
      17'd6828: data = 8'hfd;
      17'd6829: data = 8'h00;
      17'd6830: data = 8'h00;
      17'd6831: data = 8'h00;
      17'd6832: data = 8'h01;
      17'd6833: data = 8'hfd;
      17'd6834: data = 8'hfc;
      17'd6835: data = 8'h02;
      17'd6836: data = 8'h01;
      17'd6837: data = 8'hfd;
      17'd6838: data = 8'h00;
      17'd6839: data = 8'hfe;
      17'd6840: data = 8'h01;
      17'd6841: data = 8'h02;
      17'd6842: data = 8'h01;
      17'd6843: data = 8'h01;
      17'd6844: data = 8'h01;
      17'd6845: data = 8'h01;
      17'd6846: data = 8'hfe;
      17'd6847: data = 8'h00;
      17'd6848: data = 8'h02;
      17'd6849: data = 8'h04;
      17'd6850: data = 8'h00;
      17'd6851: data = 8'hfd;
      17'd6852: data = 8'h01;
      17'd6853: data = 8'h02;
      17'd6854: data = 8'h01;
      17'd6855: data = 8'h00;
      17'd6856: data = 8'h02;
      17'd6857: data = 8'h01;
      17'd6858: data = 8'h00;
      17'd6859: data = 8'hfe;
      17'd6860: data = 8'hfe;
      17'd6861: data = 8'hfe;
      17'd6862: data = 8'h00;
      17'd6863: data = 8'hfc;
      17'd6864: data = 8'hfc;
      17'd6865: data = 8'hfe;
      17'd6866: data = 8'hfd;
      17'd6867: data = 8'hfd;
      17'd6868: data = 8'hfc;
      17'd6869: data = 8'hfa;
      17'd6870: data = 8'hfc;
      17'd6871: data = 8'hfe;
      17'd6872: data = 8'h01;
      17'd6873: data = 8'hfc;
      17'd6874: data = 8'hfd;
      17'd6875: data = 8'h00;
      17'd6876: data = 8'hfa;
      17'd6877: data = 8'hfa;
      17'd6878: data = 8'hfe;
      17'd6879: data = 8'hfe;
      17'd6880: data = 8'hfc;
      17'd6881: data = 8'hfa;
      17'd6882: data = 8'hfe;
      17'd6883: data = 8'hfe;
      17'd6884: data = 8'hfc;
      17'd6885: data = 8'hfd;
      17'd6886: data = 8'hfe;
      17'd6887: data = 8'hfd;
      17'd6888: data = 8'hfd;
      17'd6889: data = 8'hfd;
      17'd6890: data = 8'hfc;
      17'd6891: data = 8'h01;
      17'd6892: data = 8'hfe;
      17'd6893: data = 8'hfc;
      17'd6894: data = 8'hfe;
      17'd6895: data = 8'hfe;
      17'd6896: data = 8'hfe;
      17'd6897: data = 8'hfd;
      17'd6898: data = 8'hfe;
      17'd6899: data = 8'hfe;
      17'd6900: data = 8'hfd;
      17'd6901: data = 8'hfa;
      17'd6902: data = 8'hfd;
      17'd6903: data = 8'h00;
      17'd6904: data = 8'hfc;
      17'd6905: data = 8'hfd;
      17'd6906: data = 8'h00;
      17'd6907: data = 8'h01;
      17'd6908: data = 8'hfd;
      17'd6909: data = 8'hfe;
      17'd6910: data = 8'hfe;
      17'd6911: data = 8'hfd;
      17'd6912: data = 8'h00;
      17'd6913: data = 8'hfe;
      17'd6914: data = 8'h01;
      17'd6915: data = 8'h02;
      17'd6916: data = 8'h01;
      17'd6917: data = 8'h01;
      17'd6918: data = 8'hfe;
      17'd6919: data = 8'hfe;
      17'd6920: data = 8'h01;
      17'd6921: data = 8'h02;
      17'd6922: data = 8'h01;
      17'd6923: data = 8'hfe;
      17'd6924: data = 8'hfd;
      17'd6925: data = 8'hfd;
      17'd6926: data = 8'h02;
      17'd6927: data = 8'h00;
      17'd6928: data = 8'h00;
      17'd6929: data = 8'h04;
      17'd6930: data = 8'h02;
      17'd6931: data = 8'hfe;
      17'd6932: data = 8'h01;
      17'd6933: data = 8'h02;
      17'd6934: data = 8'h01;
      17'd6935: data = 8'h02;
      17'd6936: data = 8'h02;
      17'd6937: data = 8'hfe;
      17'd6938: data = 8'hfe;
      17'd6939: data = 8'h01;
      17'd6940: data = 8'h01;
      17'd6941: data = 8'h01;
      17'd6942: data = 8'h04;
      17'd6943: data = 8'h01;
      17'd6944: data = 8'hfe;
      17'd6945: data = 8'h05;
      17'd6946: data = 8'h05;
      17'd6947: data = 8'h01;
      17'd6948: data = 8'hfc;
      17'd6949: data = 8'h00;
      17'd6950: data = 8'h04;
      17'd6951: data = 8'hfc;
      17'd6952: data = 8'hfc;
      17'd6953: data = 8'hfe;
      17'd6954: data = 8'hfe;
      17'd6955: data = 8'hfc;
      17'd6956: data = 8'h00;
      17'd6957: data = 8'h00;
      17'd6958: data = 8'h00;
      17'd6959: data = 8'hfe;
      17'd6960: data = 8'h00;
      17'd6961: data = 8'hfc;
      17'd6962: data = 8'hfe;
      17'd6963: data = 8'h01;
      17'd6964: data = 8'hfc;
      17'd6965: data = 8'hfd;
      17'd6966: data = 8'hfe;
      17'd6967: data = 8'hfd;
      17'd6968: data = 8'hfc;
      17'd6969: data = 8'h00;
      17'd6970: data = 8'h01;
      17'd6971: data = 8'hfd;
      17'd6972: data = 8'h00;
      17'd6973: data = 8'h01;
      17'd6974: data = 8'hfe;
      17'd6975: data = 8'h02;
      17'd6976: data = 8'h01;
      17'd6977: data = 8'hfe;
      17'd6978: data = 8'h01;
      17'd6979: data = 8'h00;
      17'd6980: data = 8'h02;
      17'd6981: data = 8'h01;
      17'd6982: data = 8'h01;
      17'd6983: data = 8'h04;
      17'd6984: data = 8'h01;
      17'd6985: data = 8'h01;
      17'd6986: data = 8'h04;
      17'd6987: data = 8'h04;
      17'd6988: data = 8'h02;
      17'd6989: data = 8'h04;
      17'd6990: data = 8'h06;
      17'd6991: data = 8'h05;
      17'd6992: data = 8'h05;
      17'd6993: data = 8'h06;
      17'd6994: data = 8'h04;
      17'd6995: data = 8'h04;
      17'd6996: data = 8'h09;
      17'd6997: data = 8'h04;
      17'd6998: data = 8'h01;
      17'd6999: data = 8'h05;
      17'd7000: data = 8'h05;
      17'd7001: data = 8'h04;
      17'd7002: data = 8'h05;
      17'd7003: data = 8'h06;
      17'd7004: data = 8'h04;
      17'd7005: data = 8'h04;
      17'd7006: data = 8'h06;
      17'd7007: data = 8'h02;
      17'd7008: data = 8'h01;
      17'd7009: data = 8'h04;
      17'd7010: data = 8'h02;
      17'd7011: data = 8'h02;
      17'd7012: data = 8'h02;
      17'd7013: data = 8'h00;
      17'd7014: data = 8'h00;
      17'd7015: data = 8'h00;
      17'd7016: data = 8'h01;
      17'd7017: data = 8'h05;
      17'd7018: data = 8'h02;
      17'd7019: data = 8'h01;
      17'd7020: data = 8'h01;
      17'd7021: data = 8'h01;
      17'd7022: data = 8'h01;
      17'd7023: data = 8'h00;
      17'd7024: data = 8'h00;
      17'd7025: data = 8'hfe;
      17'd7026: data = 8'hfe;
      17'd7027: data = 8'hfd;
      17'd7028: data = 8'hfc;
      17'd7029: data = 8'h00;
      17'd7030: data = 8'h00;
      17'd7031: data = 8'hfe;
      17'd7032: data = 8'h01;
      17'd7033: data = 8'h00;
      17'd7034: data = 8'h01;
      17'd7035: data = 8'h00;
      17'd7036: data = 8'h00;
      17'd7037: data = 8'h01;
      17'd7038: data = 8'hfd;
      17'd7039: data = 8'hfd;
      17'd7040: data = 8'hfe;
      17'd7041: data = 8'hfe;
      17'd7042: data = 8'hfe;
      17'd7043: data = 8'hfe;
      17'd7044: data = 8'hfd;
      17'd7045: data = 8'hfe;
      17'd7046: data = 8'h00;
      17'd7047: data = 8'hfe;
      17'd7048: data = 8'h00;
      17'd7049: data = 8'h00;
      17'd7050: data = 8'hfe;
      17'd7051: data = 8'hfc;
      17'd7052: data = 8'hfe;
      17'd7053: data = 8'hfe;
      17'd7054: data = 8'hfc;
      17'd7055: data = 8'hfe;
      17'd7056: data = 8'h00;
      17'd7057: data = 8'hfe;
      17'd7058: data = 8'hfc;
      17'd7059: data = 8'hfa;
      17'd7060: data = 8'hfe;
      17'd7061: data = 8'h01;
      17'd7062: data = 8'hfd;
      17'd7063: data = 8'hfc;
      17'd7064: data = 8'hfc;
      17'd7065: data = 8'h01;
      17'd7066: data = 8'h00;
      17'd7067: data = 8'hfa;
      17'd7068: data = 8'hfe;
      17'd7069: data = 8'h02;
      17'd7070: data = 8'hfd;
      17'd7071: data = 8'hfa;
      17'd7072: data = 8'hfc;
      17'd7073: data = 8'hfc;
      17'd7074: data = 8'hfd;
      17'd7075: data = 8'hfd;
      17'd7076: data = 8'hf9;
      17'd7077: data = 8'hfa;
      17'd7078: data = 8'hfa;
      17'd7079: data = 8'hf6;
      17'd7080: data = 8'hf6;
      17'd7081: data = 8'hfc;
      17'd7082: data = 8'hf6;
      17'd7083: data = 8'hf5;
      17'd7084: data = 8'hfd;
      17'd7085: data = 8'hfe;
      17'd7086: data = 8'hf9;
      17'd7087: data = 8'hfa;
      17'd7088: data = 8'hfd;
      17'd7089: data = 8'hfa;
      17'd7090: data = 8'hf9;
      17'd7091: data = 8'hfa;
      17'd7092: data = 8'hf9;
      17'd7093: data = 8'hf9;
      17'd7094: data = 8'hfc;
      17'd7095: data = 8'hfd;
      17'd7096: data = 8'hfa;
      17'd7097: data = 8'hfc;
      17'd7098: data = 8'hfe;
      17'd7099: data = 8'hfe;
      17'd7100: data = 8'h00;
      17'd7101: data = 8'h00;
      17'd7102: data = 8'hfc;
      17'd7103: data = 8'hfd;
      17'd7104: data = 8'h01;
      17'd7105: data = 8'hfe;
      17'd7106: data = 8'hfd;
      17'd7107: data = 8'hfc;
      17'd7108: data = 8'hfd;
      17'd7109: data = 8'hfe;
      17'd7110: data = 8'hfe;
      17'd7111: data = 8'h01;
      17'd7112: data = 8'h00;
      17'd7113: data = 8'h00;
      17'd7114: data = 8'h01;
      17'd7115: data = 8'h04;
      17'd7116: data = 8'h02;
      17'd7117: data = 8'hfd;
      17'd7118: data = 8'h00;
      17'd7119: data = 8'h04;
      17'd7120: data = 8'h00;
      17'd7121: data = 8'h00;
      17'd7122: data = 8'h01;
      17'd7123: data = 8'h00;
      17'd7124: data = 8'h02;
      17'd7125: data = 8'h01;
      17'd7126: data = 8'hfd;
      17'd7127: data = 8'h02;
      17'd7128: data = 8'h02;
      17'd7129: data = 8'h01;
      17'd7130: data = 8'h02;
      17'd7131: data = 8'h00;
      17'd7132: data = 8'h00;
      17'd7133: data = 8'h00;
      17'd7134: data = 8'h00;
      17'd7135: data = 8'hfd;
      17'd7136: data = 8'hfc;
      17'd7137: data = 8'hfd;
      17'd7138: data = 8'hfd;
      17'd7139: data = 8'hfc;
      17'd7140: data = 8'hfe;
      17'd7141: data = 8'hfe;
      17'd7142: data = 8'hfa;
      17'd7143: data = 8'hfc;
      17'd7144: data = 8'hfc;
      17'd7145: data = 8'hfa;
      17'd7146: data = 8'hf9;
      17'd7147: data = 8'hfa;
      17'd7148: data = 8'hf6;
      17'd7149: data = 8'hf6;
      17'd7150: data = 8'hfc;
      17'd7151: data = 8'hf9;
      17'd7152: data = 8'hf4;
      17'd7153: data = 8'hf5;
      17'd7154: data = 8'hf9;
      17'd7155: data = 8'hf9;
      17'd7156: data = 8'hf4;
      17'd7157: data = 8'hf5;
      17'd7158: data = 8'hf9;
      17'd7159: data = 8'hf4;
      17'd7160: data = 8'hf9;
      17'd7161: data = 8'hf6;
      17'd7162: data = 8'hf2;
      17'd7163: data = 8'hf4;
      17'd7164: data = 8'hf5;
      17'd7165: data = 8'hfa;
      17'd7166: data = 8'hf6;
      17'd7167: data = 8'hf4;
      17'd7168: data = 8'hf5;
      17'd7169: data = 8'hf9;
      17'd7170: data = 8'hf9;
      17'd7171: data = 8'hf9;
      17'd7172: data = 8'hf6;
      17'd7173: data = 8'hfc;
      17'd7174: data = 8'hf6;
      17'd7175: data = 8'hf5;
      17'd7176: data = 8'hfc;
      17'd7177: data = 8'hfc;
      17'd7178: data = 8'hf9;
      17'd7179: data = 8'hf6;
      17'd7180: data = 8'hfc;
      17'd7181: data = 8'hfd;
      17'd7182: data = 8'hfd;
      17'd7183: data = 8'hfc;
      17'd7184: data = 8'hfc;
      17'd7185: data = 8'hfd;
      17'd7186: data = 8'h01;
      17'd7187: data = 8'hfd;
      17'd7188: data = 8'hfc;
      17'd7189: data = 8'h01;
      17'd7190: data = 8'hfe;
      17'd7191: data = 8'hfe;
      17'd7192: data = 8'h00;
      17'd7193: data = 8'h01;
      17'd7194: data = 8'h01;
      17'd7195: data = 8'h01;
      17'd7196: data = 8'h05;
      17'd7197: data = 8'h01;
      17'd7198: data = 8'hfd;
      17'd7199: data = 8'h04;
      17'd7200: data = 8'h04;
      17'd7201: data = 8'h00;
      17'd7202: data = 8'h04;
      17'd7203: data = 8'h04;
      17'd7204: data = 8'h05;
      17'd7205: data = 8'h05;
      17'd7206: data = 8'h04;
      17'd7207: data = 8'h05;
      17'd7208: data = 8'h01;
      17'd7209: data = 8'h05;
      17'd7210: data = 8'h0a;
      17'd7211: data = 8'h00;
      17'd7212: data = 8'h04;
      17'd7213: data = 8'h05;
      17'd7214: data = 8'h02;
      17'd7215: data = 8'h0a;
      17'd7216: data = 8'h09;
      17'd7217: data = 8'h02;
      17'd7218: data = 8'h04;
      17'd7219: data = 8'h06;
      17'd7220: data = 8'h06;
      17'd7221: data = 8'h09;
      17'd7222: data = 8'h04;
      17'd7223: data = 8'h06;
      17'd7224: data = 8'h06;
      17'd7225: data = 8'h04;
      17'd7226: data = 8'h05;
      17'd7227: data = 8'h04;
      17'd7228: data = 8'h05;
      17'd7229: data = 8'h04;
      17'd7230: data = 8'h06;
      17'd7231: data = 8'h09;
      17'd7232: data = 8'h04;
      17'd7233: data = 8'h05;
      17'd7234: data = 8'h05;
      17'd7235: data = 8'h05;
      17'd7236: data = 8'h05;
      17'd7237: data = 8'h06;
      17'd7238: data = 8'h02;
      17'd7239: data = 8'h04;
      17'd7240: data = 8'h0c;
      17'd7241: data = 8'h09;
      17'd7242: data = 8'h02;
      17'd7243: data = 8'h04;
      17'd7244: data = 8'h05;
      17'd7245: data = 8'h09;
      17'd7246: data = 8'h06;
      17'd7247: data = 8'h01;
      17'd7248: data = 8'h01;
      17'd7249: data = 8'h09;
      17'd7250: data = 8'h06;
      17'd7251: data = 8'h02;
      17'd7252: data = 8'h04;
      17'd7253: data = 8'h04;
      17'd7254: data = 8'h05;
      17'd7255: data = 8'h05;
      17'd7256: data = 8'h02;
      17'd7257: data = 8'h02;
      17'd7258: data = 8'h04;
      17'd7259: data = 8'h05;
      17'd7260: data = 8'h00;
      17'd7261: data = 8'h00;
      17'd7262: data = 8'h01;
      17'd7263: data = 8'h01;
      17'd7264: data = 8'h00;
      17'd7265: data = 8'h02;
      17'd7266: data = 8'h02;
      17'd7267: data = 8'h01;
      17'd7268: data = 8'h01;
      17'd7269: data = 8'h00;
      17'd7270: data = 8'h00;
      17'd7271: data = 8'h01;
      17'd7272: data = 8'h01;
      17'd7273: data = 8'hfe;
      17'd7274: data = 8'h00;
      17'd7275: data = 8'hfe;
      17'd7276: data = 8'h00;
      17'd7277: data = 8'h01;
      17'd7278: data = 8'hfe;
      17'd7279: data = 8'h01;
      17'd7280: data = 8'h01;
      17'd7281: data = 8'h00;
      17'd7282: data = 8'hfe;
      17'd7283: data = 8'hfe;
      17'd7284: data = 8'hfe;
      17'd7285: data = 8'hfd;
      17'd7286: data = 8'hfd;
      17'd7287: data = 8'hfa;
      17'd7288: data = 8'hf9;
      17'd7289: data = 8'hfd;
      17'd7290: data = 8'hfd;
      17'd7291: data = 8'hfc;
      17'd7292: data = 8'hfa;
      17'd7293: data = 8'hfd;
      17'd7294: data = 8'hf9;
      17'd7295: data = 8'hf9;
      17'd7296: data = 8'hfc;
      17'd7297: data = 8'hf9;
      17'd7298: data = 8'hf9;
      17'd7299: data = 8'hfc;
      17'd7300: data = 8'hf9;
      17'd7301: data = 8'hf9;
      17'd7302: data = 8'hf9;
      17'd7303: data = 8'hfc;
      17'd7304: data = 8'hfa;
      17'd7305: data = 8'hf9;
      17'd7306: data = 8'hf9;
      17'd7307: data = 8'hfa;
      17'd7308: data = 8'hfd;
      17'd7309: data = 8'hfc;
      17'd7310: data = 8'hfa;
      17'd7311: data = 8'hfa;
      17'd7312: data = 8'hf9;
      17'd7313: data = 8'hfa;
      17'd7314: data = 8'hfc;
      17'd7315: data = 8'hfa;
      17'd7316: data = 8'hfa;
      17'd7317: data = 8'hfd;
      17'd7318: data = 8'hfc;
      17'd7319: data = 8'hfd;
      17'd7320: data = 8'hfd;
      17'd7321: data = 8'hfc;
      17'd7322: data = 8'hfa;
      17'd7323: data = 8'hf9;
      17'd7324: data = 8'hfa;
      17'd7325: data = 8'hfe;
      17'd7326: data = 8'hfe;
      17'd7327: data = 8'hfd;
      17'd7328: data = 8'hfd;
      17'd7329: data = 8'hfe;
      17'd7330: data = 8'h01;
      17'd7331: data = 8'h01;
      17'd7332: data = 8'hfe;
      17'd7333: data = 8'hfc;
      17'd7334: data = 8'hfe;
      17'd7335: data = 8'h01;
      17'd7336: data = 8'hfc;
      17'd7337: data = 8'hf6;
      17'd7338: data = 8'hfd;
      17'd7339: data = 8'h00;
      17'd7340: data = 8'hfe;
      17'd7341: data = 8'hfe;
      17'd7342: data = 8'hfc;
      17'd7343: data = 8'hfe;
      17'd7344: data = 8'h01;
      17'd7345: data = 8'hfd;
      17'd7346: data = 8'hfe;
      17'd7347: data = 8'h01;
      17'd7348: data = 8'hfc;
      17'd7349: data = 8'hfa;
      17'd7350: data = 8'hfd;
      17'd7351: data = 8'hfa;
      17'd7352: data = 8'hf9;
      17'd7353: data = 8'hfc;
      17'd7354: data = 8'hfc;
      17'd7355: data = 8'hfa;
      17'd7356: data = 8'hfc;
      17'd7357: data = 8'hfc;
      17'd7358: data = 8'hf9;
      17'd7359: data = 8'hfc;
      17'd7360: data = 8'hfd;
      17'd7361: data = 8'hf9;
      17'd7362: data = 8'hfa;
      17'd7363: data = 8'hfc;
      17'd7364: data = 8'hfc;
      17'd7365: data = 8'hfc;
      17'd7366: data = 8'hf9;
      17'd7367: data = 8'hf5;
      17'd7368: data = 8'hf9;
      17'd7369: data = 8'hfd;
      17'd7370: data = 8'hfc;
      17'd7371: data = 8'hf5;
      17'd7372: data = 8'hf9;
      17'd7373: data = 8'hfe;
      17'd7374: data = 8'hfa;
      17'd7375: data = 8'hfc;
      17'd7376: data = 8'hfc;
      17'd7377: data = 8'hfd;
      17'd7378: data = 8'hfd;
      17'd7379: data = 8'hfc;
      17'd7380: data = 8'hfd;
      17'd7381: data = 8'hfd;
      17'd7382: data = 8'hfc;
      17'd7383: data = 8'h00;
      17'd7384: data = 8'hfe;
      17'd7385: data = 8'hfc;
      17'd7386: data = 8'hfe;
      17'd7387: data = 8'hfa;
      17'd7388: data = 8'hfc;
      17'd7389: data = 8'h00;
      17'd7390: data = 8'h00;
      17'd7391: data = 8'hfe;
      17'd7392: data = 8'h00;
      17'd7393: data = 8'h01;
      17'd7394: data = 8'hfe;
      17'd7395: data = 8'hfd;
      17'd7396: data = 8'h00;
      17'd7397: data = 8'h01;
      17'd7398: data = 8'h00;
      17'd7399: data = 8'h00;
      17'd7400: data = 8'hfe;
      17'd7401: data = 8'hfe;
      17'd7402: data = 8'h01;
      17'd7403: data = 8'h01;
      17'd7404: data = 8'h00;
      17'd7405: data = 8'h04;
      17'd7406: data = 8'h02;
      17'd7407: data = 8'h02;
      17'd7408: data = 8'h04;
      17'd7409: data = 8'h04;
      17'd7410: data = 8'h02;
      17'd7411: data = 8'h02;
      17'd7412: data = 8'h02;
      17'd7413: data = 8'h04;
      17'd7414: data = 8'h02;
      17'd7415: data = 8'h01;
      17'd7416: data = 8'h02;
      17'd7417: data = 8'h05;
      17'd7418: data = 8'h05;
      17'd7419: data = 8'h05;
      17'd7420: data = 8'h05;
      17'd7421: data = 8'h02;
      17'd7422: data = 8'h02;
      17'd7423: data = 8'h05;
      17'd7424: data = 8'h01;
      17'd7425: data = 8'h02;
      17'd7426: data = 8'h05;
      17'd7427: data = 8'h01;
      17'd7428: data = 8'h05;
      17'd7429: data = 8'h02;
      17'd7430: data = 8'h00;
      17'd7431: data = 8'h02;
      17'd7432: data = 8'h04;
      17'd7433: data = 8'h04;
      17'd7434: data = 8'h02;
      17'd7435: data = 8'h02;
      17'd7436: data = 8'h02;
      17'd7437: data = 8'h00;
      17'd7438: data = 8'h04;
      17'd7439: data = 8'h04;
      17'd7440: data = 8'hfe;
      17'd7441: data = 8'h02;
      17'd7442: data = 8'h01;
      17'd7443: data = 8'h01;
      17'd7444: data = 8'h02;
      17'd7445: data = 8'h00;
      17'd7446: data = 8'h02;
      17'd7447: data = 8'h02;
      17'd7448: data = 8'h01;
      17'd7449: data = 8'h01;
      17'd7450: data = 8'h01;
      17'd7451: data = 8'h05;
      17'd7452: data = 8'h05;
      17'd7453: data = 8'h02;
      17'd7454: data = 8'h02;
      17'd7455: data = 8'h02;
      17'd7456: data = 8'h02;
      17'd7457: data = 8'h04;
      17'd7458: data = 8'h05;
      17'd7459: data = 8'h02;
      17'd7460: data = 8'h02;
      17'd7461: data = 8'h04;
      17'd7462: data = 8'h04;
      17'd7463: data = 8'h04;
      17'd7464: data = 8'h05;
      17'd7465: data = 8'h02;
      17'd7466: data = 8'h00;
      17'd7467: data = 8'h05;
      17'd7468: data = 8'h05;
      17'd7469: data = 8'h04;
      17'd7470: data = 8'h04;
      17'd7471: data = 8'h01;
      17'd7472: data = 8'h02;
      17'd7473: data = 8'h05;
      17'd7474: data = 8'h04;
      17'd7475: data = 8'h01;
      17'd7476: data = 8'h01;
      17'd7477: data = 8'h05;
      17'd7478: data = 8'h06;
      17'd7479: data = 8'h02;
      17'd7480: data = 8'h02;
      17'd7481: data = 8'h05;
      17'd7482: data = 8'h04;
      17'd7483: data = 8'h02;
      17'd7484: data = 8'h01;
      17'd7485: data = 8'h02;
      17'd7486: data = 8'h05;
      17'd7487: data = 8'h04;
      17'd7488: data = 8'h02;
      17'd7489: data = 8'h01;
      17'd7490: data = 8'h01;
      17'd7491: data = 8'h02;
      17'd7492: data = 8'h01;
      17'd7493: data = 8'h04;
      17'd7494: data = 8'h05;
      17'd7495: data = 8'h01;
      17'd7496: data = 8'hfe;
      17'd7497: data = 8'h02;
      17'd7498: data = 8'h02;
      17'd7499: data = 8'h01;
      17'd7500: data = 8'hfe;
      17'd7501: data = 8'hfe;
      17'd7502: data = 8'h02;
      17'd7503: data = 8'h01;
      17'd7504: data = 8'hfd;
      17'd7505: data = 8'hfe;
      17'd7506: data = 8'h00;
      17'd7507: data = 8'h01;
      17'd7508: data = 8'hfe;
      17'd7509: data = 8'hfc;
      17'd7510: data = 8'hfd;
      17'd7511: data = 8'h01;
      17'd7512: data = 8'h00;
      17'd7513: data = 8'hfe;
      17'd7514: data = 8'hfc;
      17'd7515: data = 8'hfd;
      17'd7516: data = 8'h01;
      17'd7517: data = 8'h02;
      17'd7518: data = 8'hfe;
      17'd7519: data = 8'hfd;
      17'd7520: data = 8'h00;
      17'd7521: data = 8'h01;
      17'd7522: data = 8'h01;
      17'd7523: data = 8'h00;
      17'd7524: data = 8'h01;
      17'd7525: data = 8'h00;
      17'd7526: data = 8'h00;
      17'd7527: data = 8'h01;
      17'd7528: data = 8'h02;
      17'd7529: data = 8'h01;
      17'd7530: data = 8'h00;
      17'd7531: data = 8'hfe;
      17'd7532: data = 8'h00;
      17'd7533: data = 8'h00;
      17'd7534: data = 8'h01;
      17'd7535: data = 8'h02;
      17'd7536: data = 8'h01;
      17'd7537: data = 8'h01;
      17'd7538: data = 8'h02;
      17'd7539: data = 8'h04;
      17'd7540: data = 8'h01;
      17'd7541: data = 8'h01;
      17'd7542: data = 8'h02;
      17'd7543: data = 8'h02;
      17'd7544: data = 8'h00;
      17'd7545: data = 8'h02;
      17'd7546: data = 8'h02;
      17'd7547: data = 8'hfe;
      17'd7548: data = 8'h00;
      17'd7549: data = 8'h02;
      17'd7550: data = 8'h02;
      17'd7551: data = 8'h00;
      17'd7552: data = 8'h00;
      17'd7553: data = 8'h00;
      17'd7554: data = 8'h02;
      17'd7555: data = 8'h02;
      17'd7556: data = 8'h00;
      17'd7557: data = 8'h00;
      17'd7558: data = 8'h01;
      17'd7559: data = 8'h01;
      17'd7560: data = 8'h00;
      17'd7561: data = 8'hfd;
      17'd7562: data = 8'hfd;
      17'd7563: data = 8'hfe;
      17'd7564: data = 8'hfd;
      17'd7565: data = 8'h00;
      17'd7566: data = 8'h00;
      17'd7567: data = 8'hfe;
      17'd7568: data = 8'hfd;
      17'd7569: data = 8'h00;
      17'd7570: data = 8'h00;
      17'd7571: data = 8'hfa;
      17'd7572: data = 8'hfd;
      17'd7573: data = 8'hfe;
      17'd7574: data = 8'hfc;
      17'd7575: data = 8'hfc;
      17'd7576: data = 8'hf9;
      17'd7577: data = 8'hfa;
      17'd7578: data = 8'hfd;
      17'd7579: data = 8'hfa;
      17'd7580: data = 8'hf6;
      17'd7581: data = 8'hfa;
      17'd7582: data = 8'hfa;
      17'd7583: data = 8'hfe;
      17'd7584: data = 8'hfd;
      17'd7585: data = 8'hf9;
      17'd7586: data = 8'hfc;
      17'd7587: data = 8'hfc;
      17'd7588: data = 8'hf9;
      17'd7589: data = 8'hfa;
      17'd7590: data = 8'hf9;
      17'd7591: data = 8'hf6;
      17'd7592: data = 8'hfa;
      17'd7593: data = 8'hfc;
      17'd7594: data = 8'hfc;
      17'd7595: data = 8'hfa;
      17'd7596: data = 8'hfc;
      17'd7597: data = 8'hfe;
      17'd7598: data = 8'hfe;
      17'd7599: data = 8'hfd;
      17'd7600: data = 8'hfd;
      17'd7601: data = 8'hfc;
      17'd7602: data = 8'hfc;
      17'd7603: data = 8'hfd;
      17'd7604: data = 8'hfd;
      17'd7605: data = 8'hfc;
      17'd7606: data = 8'hfa;
      17'd7607: data = 8'hfa;
      17'd7608: data = 8'hfa;
      17'd7609: data = 8'hfc;
      17'd7610: data = 8'hfd;
      17'd7611: data = 8'hfc;
      17'd7612: data = 8'hfe;
      17'd7613: data = 8'h01;
      17'd7614: data = 8'h01;
      17'd7615: data = 8'hfd;
      17'd7616: data = 8'hfd;
      17'd7617: data = 8'h00;
      17'd7618: data = 8'h00;
      17'd7619: data = 8'h00;
      17'd7620: data = 8'h00;
      17'd7621: data = 8'hfd;
      17'd7622: data = 8'hfe;
      17'd7623: data = 8'h02;
      17'd7624: data = 8'h00;
      17'd7625: data = 8'hfd;
      17'd7626: data = 8'h00;
      17'd7627: data = 8'h02;
      17'd7628: data = 8'h00;
      17'd7629: data = 8'h02;
      17'd7630: data = 8'h00;
      17'd7631: data = 8'h00;
      17'd7632: data = 8'h02;
      17'd7633: data = 8'h00;
      17'd7634: data = 8'hfe;
      17'd7635: data = 8'h02;
      17'd7636: data = 8'h02;
      17'd7637: data = 8'h00;
      17'd7638: data = 8'h00;
      17'd7639: data = 8'h01;
      17'd7640: data = 8'h00;
      17'd7641: data = 8'hfe;
      17'd7642: data = 8'h00;
      17'd7643: data = 8'h00;
      17'd7644: data = 8'h00;
      17'd7645: data = 8'hfe;
      17'd7646: data = 8'hfd;
      17'd7647: data = 8'hfe;
      17'd7648: data = 8'h00;
      17'd7649: data = 8'h01;
      17'd7650: data = 8'hfd;
      17'd7651: data = 8'hfa;
      17'd7652: data = 8'hfd;
      17'd7653: data = 8'hfd;
      17'd7654: data = 8'hfd;
      17'd7655: data = 8'hfe;
      17'd7656: data = 8'hfe;
      17'd7657: data = 8'hfc;
      17'd7658: data = 8'hfc;
      17'd7659: data = 8'h00;
      17'd7660: data = 8'hfd;
      17'd7661: data = 8'hfa;
      17'd7662: data = 8'hfc;
      17'd7663: data = 8'hfd;
      17'd7664: data = 8'hfd;
      17'd7665: data = 8'hfa;
      17'd7666: data = 8'hfc;
      17'd7667: data = 8'h00;
      17'd7668: data = 8'hfd;
      17'd7669: data = 8'hf9;
      17'd7670: data = 8'hfc;
      17'd7671: data = 8'hfe;
      17'd7672: data = 8'hfd;
      17'd7673: data = 8'hfc;
      17'd7674: data = 8'hfa;
      17'd7675: data = 8'hfd;
      17'd7676: data = 8'hfd;
      17'd7677: data = 8'hfc;
      17'd7678: data = 8'hfc;
      17'd7679: data = 8'hfc;
      17'd7680: data = 8'hfa;
      17'd7681: data = 8'hfc;
      17'd7682: data = 8'hfd;
      17'd7683: data = 8'hfc;
      17'd7684: data = 8'hfd;
      17'd7685: data = 8'h00;
      17'd7686: data = 8'hfd;
      17'd7687: data = 8'hfc;
      17'd7688: data = 8'hfe;
      17'd7689: data = 8'hfe;
      17'd7690: data = 8'hfe;
      17'd7691: data = 8'hfe;
      17'd7692: data = 8'hfd;
      17'd7693: data = 8'hfd;
      17'd7694: data = 8'h00;
      17'd7695: data = 8'hfe;
      17'd7696: data = 8'hfc;
      17'd7697: data = 8'h01;
      17'd7698: data = 8'h01;
      17'd7699: data = 8'hfd;
      17'd7700: data = 8'hfd;
      17'd7701: data = 8'h01;
      17'd7702: data = 8'h00;
      17'd7703: data = 8'hfe;
      17'd7704: data = 8'h00;
      17'd7705: data = 8'hfe;
      17'd7706: data = 8'hfd;
      17'd7707: data = 8'h00;
      17'd7708: data = 8'h01;
      17'd7709: data = 8'h02;
      17'd7710: data = 8'h04;
      17'd7711: data = 8'h00;
      17'd7712: data = 8'h00;
      17'd7713: data = 8'h01;
      17'd7714: data = 8'h01;
      17'd7715: data = 8'hfd;
      17'd7716: data = 8'hfd;
      17'd7717: data = 8'h00;
      17'd7718: data = 8'h00;
      17'd7719: data = 8'h00;
      17'd7720: data = 8'h00;
      17'd7721: data = 8'h00;
      17'd7722: data = 8'hfd;
      17'd7723: data = 8'h01;
      17'd7724: data = 8'h04;
      17'd7725: data = 8'h04;
      17'd7726: data = 8'h02;
      17'd7727: data = 8'h00;
      17'd7728: data = 8'h00;
      17'd7729: data = 8'h01;
      17'd7730: data = 8'h02;
      17'd7731: data = 8'h01;
      17'd7732: data = 8'h01;
      17'd7733: data = 8'h01;
      17'd7734: data = 8'h04;
      17'd7735: data = 8'h05;
      17'd7736: data = 8'h04;
      17'd7737: data = 8'h04;
      17'd7738: data = 8'h06;
      17'd7739: data = 8'h05;
      17'd7740: data = 8'h05;
      17'd7741: data = 8'h05;
      17'd7742: data = 8'h02;
      17'd7743: data = 8'h02;
      17'd7744: data = 8'h05;
      17'd7745: data = 8'h04;
      17'd7746: data = 8'h04;
      17'd7747: data = 8'h06;
      17'd7748: data = 8'h02;
      17'd7749: data = 8'h02;
      17'd7750: data = 8'h05;
      17'd7751: data = 8'h06;
      17'd7752: data = 8'h05;
      17'd7753: data = 8'h05;
      17'd7754: data = 8'h02;
      17'd7755: data = 8'h05;
      17'd7756: data = 8'h06;
      17'd7757: data = 8'h01;
      17'd7758: data = 8'h02;
      17'd7759: data = 8'h01;
      17'd7760: data = 8'h01;
      17'd7761: data = 8'h02;
      17'd7762: data = 8'h02;
      17'd7763: data = 8'h00;
      17'd7764: data = 8'h00;
      17'd7765: data = 8'h04;
      17'd7766: data = 8'h01;
      17'd7767: data = 8'hfe;
      17'd7768: data = 8'h00;
      17'd7769: data = 8'h00;
      17'd7770: data = 8'h04;
      17'd7771: data = 8'h02;
      17'd7772: data = 8'hfd;
      17'd7773: data = 8'hfe;
      17'd7774: data = 8'h01;
      17'd7775: data = 8'h00;
      17'd7776: data = 8'hfe;
      17'd7777: data = 8'h01;
      17'd7778: data = 8'h00;
      17'd7779: data = 8'hfa;
      17'd7780: data = 8'h00;
      17'd7781: data = 8'h02;
      17'd7782: data = 8'hfe;
      17'd7783: data = 8'hfe;
      17'd7784: data = 8'h00;
      17'd7785: data = 8'h01;
      17'd7786: data = 8'h00;
      17'd7787: data = 8'hfe;
      17'd7788: data = 8'hfd;
      17'd7789: data = 8'hfe;
      17'd7790: data = 8'h00;
      17'd7791: data = 8'h00;
      17'd7792: data = 8'hfd;
      17'd7793: data = 8'h00;
      17'd7794: data = 8'h00;
      17'd7795: data = 8'hfe;
      17'd7796: data = 8'h01;
      17'd7797: data = 8'hfd;
      17'd7798: data = 8'hfd;
      17'd7799: data = 8'hfe;
      17'd7800: data = 8'h00;
      17'd7801: data = 8'h01;
      17'd7802: data = 8'hfe;
      17'd7803: data = 8'hfe;
      17'd7804: data = 8'h00;
      17'd7805: data = 8'h02;
      17'd7806: data = 8'h00;
      17'd7807: data = 8'hfe;
      17'd7808: data = 8'h00;
      17'd7809: data = 8'h00;
      17'd7810: data = 8'h00;
      17'd7811: data = 8'h00;
      17'd7812: data = 8'hfd;
      17'd7813: data = 8'hfd;
      17'd7814: data = 8'h00;
      17'd7815: data = 8'h01;
      17'd7816: data = 8'hfe;
      17'd7817: data = 8'hfe;
      17'd7818: data = 8'h01;
      17'd7819: data = 8'h01;
      17'd7820: data = 8'h01;
      17'd7821: data = 8'hfe;
      17'd7822: data = 8'hfe;
      17'd7823: data = 8'h00;
      17'd7824: data = 8'h00;
      17'd7825: data = 8'h00;
      17'd7826: data = 8'hfd;
      17'd7827: data = 8'hfc;
      17'd7828: data = 8'hfd;
      17'd7829: data = 8'hfe;
      17'd7830: data = 8'hfd;
      17'd7831: data = 8'hfc;
      17'd7832: data = 8'hfe;
      17'd7833: data = 8'hfd;
      17'd7834: data = 8'hfd;
      17'd7835: data = 8'hfe;
      17'd7836: data = 8'hfe;
      17'd7837: data = 8'h01;
      17'd7838: data = 8'hfe;
      17'd7839: data = 8'hfc;
      17'd7840: data = 8'hfe;
      17'd7841: data = 8'hfe;
      17'd7842: data = 8'hfd;
      17'd7843: data = 8'hfe;
      17'd7844: data = 8'hfe;
      17'd7845: data = 8'hfc;
      17'd7846: data = 8'hfd;
      17'd7847: data = 8'hfd;
      17'd7848: data = 8'hfe;
      17'd7849: data = 8'hfe;
      17'd7850: data = 8'h01;
      17'd7851: data = 8'hfd;
      17'd7852: data = 8'hfc;
      17'd7853: data = 8'h00;
      17'd7854: data = 8'h00;
      17'd7855: data = 8'hfc;
      17'd7856: data = 8'hfc;
      17'd7857: data = 8'hfd;
      17'd7858: data = 8'hfa;
      17'd7859: data = 8'hfd;
      17'd7860: data = 8'hfe;
      17'd7861: data = 8'hfc;
      17'd7862: data = 8'hfd;
      17'd7863: data = 8'hfc;
      17'd7864: data = 8'hfc;
      17'd7865: data = 8'hfd;
      17'd7866: data = 8'hfe;
      17'd7867: data = 8'h01;
      17'd7868: data = 8'h00;
      17'd7869: data = 8'hfc;
      17'd7870: data = 8'hfd;
      17'd7871: data = 8'hfe;
      17'd7872: data = 8'hfc;
      17'd7873: data = 8'hfd;
      17'd7874: data = 8'hfe;
      17'd7875: data = 8'hfd;
      17'd7876: data = 8'hfe;
      17'd7877: data = 8'hfd;
      17'd7878: data = 8'hfd;
      17'd7879: data = 8'h00;
      17'd7880: data = 8'h01;
      17'd7881: data = 8'hfe;
      17'd7882: data = 8'hfd;
      17'd7883: data = 8'h00;
      17'd7884: data = 8'h00;
      17'd7885: data = 8'hfd;
      17'd7886: data = 8'hfd;
      17'd7887: data = 8'h00;
      17'd7888: data = 8'hfd;
      17'd7889: data = 8'hfd;
      17'd7890: data = 8'hfd;
      17'd7891: data = 8'hfc;
      17'd7892: data = 8'hfe;
      17'd7893: data = 8'hfd;
      17'd7894: data = 8'hfc;
      17'd7895: data = 8'hfe;
      17'd7896: data = 8'h00;
      17'd7897: data = 8'hfe;
      17'd7898: data = 8'hfd;
      17'd7899: data = 8'h00;
      17'd7900: data = 8'hfd;
      17'd7901: data = 8'hfe;
      17'd7902: data = 8'h00;
      17'd7903: data = 8'h01;
      17'd7904: data = 8'h00;
      17'd7905: data = 8'h00;
      17'd7906: data = 8'h00;
      17'd7907: data = 8'h01;
      17'd7908: data = 8'h00;
      17'd7909: data = 8'hfe;
      17'd7910: data = 8'hfe;
      17'd7911: data = 8'hfd;
      17'd7912: data = 8'h00;
      17'd7913: data = 8'hfe;
      17'd7914: data = 8'h00;
      17'd7915: data = 8'h00;
      17'd7916: data = 8'h00;
      17'd7917: data = 8'h02;
      17'd7918: data = 8'hfd;
      17'd7919: data = 8'hfd;
      17'd7920: data = 8'h00;
      17'd7921: data = 8'hfe;
      17'd7922: data = 8'hfe;
      17'd7923: data = 8'h00;
      17'd7924: data = 8'hfe;
      17'd7925: data = 8'hfa;
      17'd7926: data = 8'hfa;
      17'd7927: data = 8'hfd;
      17'd7928: data = 8'hfc;
      17'd7929: data = 8'hfd;
      17'd7930: data = 8'h00;
      17'd7931: data = 8'hfc;
      17'd7932: data = 8'hfd;
      17'd7933: data = 8'h01;
      17'd7934: data = 8'h00;
      17'd7935: data = 8'hfd;
      17'd7936: data = 8'hfd;
      17'd7937: data = 8'h00;
      17'd7938: data = 8'hfe;
      17'd7939: data = 8'hfc;
      17'd7940: data = 8'h00;
      17'd7941: data = 8'h00;
      17'd7942: data = 8'hfc;
      17'd7943: data = 8'hfd;
      17'd7944: data = 8'h01;
      17'd7945: data = 8'h00;
      17'd7946: data = 8'h00;
      17'd7947: data = 8'h02;
      17'd7948: data = 8'h01;
      17'd7949: data = 8'h00;
      17'd7950: data = 8'h04;
      17'd7951: data = 8'h04;
      17'd7952: data = 8'h01;
      17'd7953: data = 8'h04;
      17'd7954: data = 8'h04;
      17'd7955: data = 8'h00;
      17'd7956: data = 8'hfe;
      17'd7957: data = 8'h02;
      17'd7958: data = 8'h00;
      17'd7959: data = 8'h01;
      17'd7960: data = 8'h04;
      17'd7961: data = 8'h01;
      17'd7962: data = 8'hfe;
      17'd7963: data = 8'h02;
      17'd7964: data = 8'h05;
      17'd7965: data = 8'h00;
      17'd7966: data = 8'h02;
      17'd7967: data = 8'h02;
      17'd7968: data = 8'h01;
      17'd7969: data = 8'h01;
      17'd7970: data = 8'h00;
      17'd7971: data = 8'h01;
      17'd7972: data = 8'h00;
      17'd7973: data = 8'h01;
      17'd7974: data = 8'h01;
      17'd7975: data = 8'h00;
      17'd7976: data = 8'h02;
      17'd7977: data = 8'hfe;
      17'd7978: data = 8'hfe;
      17'd7979: data = 8'h00;
      17'd7980: data = 8'h00;
      17'd7981: data = 8'hfe;
      17'd7982: data = 8'hfa;
      17'd7983: data = 8'h00;
      17'd7984: data = 8'h01;
      17'd7985: data = 8'hfe;
      17'd7986: data = 8'hfd;
      17'd7987: data = 8'hfe;
      17'd7988: data = 8'h00;
      17'd7989: data = 8'hfe;
      17'd7990: data = 8'h01;
      17'd7991: data = 8'h00;
      17'd7992: data = 8'hfd;
      17'd7993: data = 8'hfe;
      17'd7994: data = 8'h00;
      17'd7995: data = 8'hfd;
      17'd7996: data = 8'hfe;
      17'd7997: data = 8'h00;
      17'd7998: data = 8'hfe;
      17'd7999: data = 8'h00;
      17'd8000: data = 8'h02;
      17'd8001: data = 8'h01;
      17'd8002: data = 8'h01;
      17'd8003: data = 8'h00;
      17'd8004: data = 8'h02;
      17'd8005: data = 8'h02;
      17'd8006: data = 8'hfc;
      17'd8007: data = 8'hfe;
      17'd8008: data = 8'h02;
      17'd8009: data = 8'h01;
      17'd8010: data = 8'hfe;
      17'd8011: data = 8'h01;
      17'd8012: data = 8'h01;
      17'd8013: data = 8'h01;
      17'd8014: data = 8'h01;
      17'd8015: data = 8'h00;
      17'd8016: data = 8'h01;
      17'd8017: data = 8'h04;
      17'd8018: data = 8'h02;
      17'd8019: data = 8'h00;
      17'd8020: data = 8'h01;
      17'd8021: data = 8'h02;
      17'd8022: data = 8'hfe;
      17'd8023: data = 8'hfd;
      17'd8024: data = 8'h00;
      17'd8025: data = 8'h00;
      17'd8026: data = 8'hfe;
      17'd8027: data = 8'h01;
      17'd8028: data = 8'h02;
      17'd8029: data = 8'h01;
      17'd8030: data = 8'h02;
      17'd8031: data = 8'h01;
      17'd8032: data = 8'hfe;
      17'd8033: data = 8'h01;
      17'd8034: data = 8'h00;
      17'd8035: data = 8'hfe;
      17'd8036: data = 8'h00;
      17'd8037: data = 8'h00;
      17'd8038: data = 8'h00;
      17'd8039: data = 8'h00;
      17'd8040: data = 8'hfe;
      17'd8041: data = 8'hfd;
      17'd8042: data = 8'hfd;
      17'd8043: data = 8'hfe;
      17'd8044: data = 8'h00;
      17'd8045: data = 8'h01;
      17'd8046: data = 8'h01;
      17'd8047: data = 8'h01;
      17'd8048: data = 8'hfe;
      17'd8049: data = 8'hfc;
      17'd8050: data = 8'hfd;
      17'd8051: data = 8'hfe;
      17'd8052: data = 8'hfe;
      17'd8053: data = 8'hfd;
      17'd8054: data = 8'hfd;
      17'd8055: data = 8'hfd;
      17'd8056: data = 8'hfd;
      17'd8057: data = 8'h00;
      17'd8058: data = 8'hfe;
      17'd8059: data = 8'hfd;
      17'd8060: data = 8'h00;
      17'd8061: data = 8'h00;
      17'd8062: data = 8'hfd;
      17'd8063: data = 8'hfd;
      17'd8064: data = 8'hfe;
      17'd8065: data = 8'h00;
      17'd8066: data = 8'hfe;
      17'd8067: data = 8'h00;
      17'd8068: data = 8'hfe;
      17'd8069: data = 8'hfa;
      17'd8070: data = 8'hfc;
      17'd8071: data = 8'hfd;
      17'd8072: data = 8'hfc;
      17'd8073: data = 8'hfe;
      17'd8074: data = 8'hfe;
      17'd8075: data = 8'hfd;
      17'd8076: data = 8'hfe;
      17'd8077: data = 8'h00;
      17'd8078: data = 8'hfd;
      17'd8079: data = 8'hfd;
      17'd8080: data = 8'hfe;
      17'd8081: data = 8'hfd;
      17'd8082: data = 8'hfe;
      17'd8083: data = 8'h00;
      17'd8084: data = 8'hfd;
      17'd8085: data = 8'hfd;
      17'd8086: data = 8'hfc;
      17'd8087: data = 8'h01;
      17'd8088: data = 8'h01;
      17'd8089: data = 8'hfc;
      17'd8090: data = 8'hfd;
      17'd8091: data = 8'hfe;
      17'd8092: data = 8'h00;
      17'd8093: data = 8'h00;
      17'd8094: data = 8'hfe;
      17'd8095: data = 8'h00;
      17'd8096: data = 8'h00;
      17'd8097: data = 8'hfe;
      17'd8098: data = 8'h01;
      17'd8099: data = 8'h02;
      17'd8100: data = 8'h01;
      17'd8101: data = 8'hfe;
      17'd8102: data = 8'hfe;
      17'd8103: data = 8'h00;
      17'd8104: data = 8'hfe;
      17'd8105: data = 8'hfd;
      17'd8106: data = 8'hfe;
      17'd8107: data = 8'h00;
      17'd8108: data = 8'h00;
      17'd8109: data = 8'h00;
      17'd8110: data = 8'h01;
      17'd8111: data = 8'h01;
      17'd8112: data = 8'h00;
      17'd8113: data = 8'h01;
      17'd8114: data = 8'h01;
      17'd8115: data = 8'hfe;
      17'd8116: data = 8'hfd;
      17'd8117: data = 8'hfe;
      17'd8118: data = 8'hfe;
      17'd8119: data = 8'hfe;
      17'd8120: data = 8'hfe;
      17'd8121: data = 8'hfe;
      17'd8122: data = 8'hfe;
      17'd8123: data = 8'hfc;
      17'd8124: data = 8'h00;
      17'd8125: data = 8'h01;
      17'd8126: data = 8'hfd;
      17'd8127: data = 8'hfd;
      17'd8128: data = 8'h01;
      17'd8129: data = 8'h01;
      17'd8130: data = 8'hfd;
      17'd8131: data = 8'hfd;
      17'd8132: data = 8'hfd;
      17'd8133: data = 8'hfd;
      17'd8134: data = 8'hfe;
      17'd8135: data = 8'hfe;
      17'd8136: data = 8'hfe;
      17'd8137: data = 8'h00;
      17'd8138: data = 8'hfe;
      17'd8139: data = 8'hfd;
      17'd8140: data = 8'hfd;
      17'd8141: data = 8'h00;
      17'd8142: data = 8'h00;
      17'd8143: data = 8'hfd;
      17'd8144: data = 8'hfc;
      17'd8145: data = 8'hfd;
      17'd8146: data = 8'hfc;
      17'd8147: data = 8'hfc;
      17'd8148: data = 8'hfd;
      17'd8149: data = 8'hfe;
      17'd8150: data = 8'hfe;
      17'd8151: data = 8'h00;
      17'd8152: data = 8'hfe;
      17'd8153: data = 8'hfd;
      17'd8154: data = 8'hfd;
      17'd8155: data = 8'hfc;
      17'd8156: data = 8'hfd;
      17'd8157: data = 8'hfe;
      17'd8158: data = 8'h00;
      17'd8159: data = 8'h04;
      17'd8160: data = 8'hf6;
      17'd8161: data = 8'h02;
      17'd8162: data = 8'h0c;
      17'd8163: data = 8'h00;
      17'd8164: data = 8'h02;
      17'd8165: data = 8'hfe;
      17'd8166: data = 8'hfd;
      17'd8167: data = 8'h06;
      17'd8168: data = 8'h02;
      17'd8169: data = 8'h02;
      17'd8170: data = 8'h06;
      17'd8171: data = 8'h00;
      17'd8172: data = 8'h00;
      17'd8173: data = 8'h04;
      17'd8174: data = 8'h02;
      17'd8175: data = 8'h02;
      17'd8176: data = 8'h01;
      17'd8177: data = 8'h01;
      17'd8178: data = 8'h04;
      17'd8179: data = 8'h04;
      17'd8180: data = 8'h06;
      17'd8181: data = 8'h02;
      17'd8182: data = 8'hf2;
      17'd8183: data = 8'hf9;
      17'd8184: data = 8'h04;
      17'd8185: data = 8'h00;
      17'd8186: data = 8'h00;
      17'd8187: data = 8'h02;
      17'd8188: data = 8'h01;
      17'd8189: data = 8'h05;
      17'd8190: data = 8'h00;
      17'd8191: data = 8'hfe;
      17'd8192: data = 8'h05;
      17'd8193: data = 8'h01;
      17'd8194: data = 8'hfd;
      17'd8195: data = 8'hfd;
      17'd8196: data = 8'hfe;
      17'd8197: data = 8'h01;
      17'd8198: data = 8'hfd;
      17'd8199: data = 8'hf6;
      17'd8200: data = 8'hfc;
      17'd8201: data = 8'hfe;
      17'd8202: data = 8'h01;
      17'd8203: data = 8'h04;
      17'd8204: data = 8'hfe;
      17'd8205: data = 8'hfc;
      17'd8206: data = 8'hfe;
      17'd8207: data = 8'h00;
      17'd8208: data = 8'h04;
      17'd8209: data = 8'h02;
      17'd8210: data = 8'h00;
      17'd8211: data = 8'h02;
      17'd8212: data = 8'hfe;
      17'd8213: data = 8'hfe;
      17'd8214: data = 8'h00;
      17'd8215: data = 8'h00;
      17'd8216: data = 8'hfd;
      17'd8217: data = 8'hfd;
      17'd8218: data = 8'h00;
      17'd8219: data = 8'h00;
      17'd8220: data = 8'h00;
      17'd8221: data = 8'hfe;
      17'd8222: data = 8'h00;
      17'd8223: data = 8'h01;
      17'd8224: data = 8'h00;
      17'd8225: data = 8'hfd;
      17'd8226: data = 8'h00;
      17'd8227: data = 8'hfd;
      17'd8228: data = 8'h00;
      17'd8229: data = 8'hfd;
      17'd8230: data = 8'hfc;
      17'd8231: data = 8'h01;
      17'd8232: data = 8'h01;
      17'd8233: data = 8'h00;
      17'd8234: data = 8'h01;
      17'd8235: data = 8'h01;
      17'd8236: data = 8'h00;
      17'd8237: data = 8'h02;
      17'd8238: data = 8'h01;
      17'd8239: data = 8'h00;
      17'd8240: data = 8'hfa;
      17'd8241: data = 8'h00;
      17'd8242: data = 8'h00;
      17'd8243: data = 8'h05;
      17'd8244: data = 8'h00;
      17'd8245: data = 8'hf6;
      17'd8246: data = 8'h01;
      17'd8247: data = 8'h00;
      17'd8248: data = 8'h00;
      17'd8249: data = 8'h01;
      17'd8250: data = 8'h00;
      17'd8251: data = 8'h02;
      17'd8252: data = 8'h01;
      17'd8253: data = 8'h00;
      17'd8254: data = 8'h04;
      17'd8255: data = 8'hfd;
      17'd8256: data = 8'hfa;
      17'd8257: data = 8'hfa;
      17'd8258: data = 8'hf9;
      17'd8259: data = 8'hfd;
      17'd8260: data = 8'hfc;
      17'd8261: data = 8'hfe;
      17'd8262: data = 8'hfd;
      17'd8263: data = 8'hfe;
      17'd8264: data = 8'h01;
      17'd8265: data = 8'h00;
      17'd8266: data = 8'hfc;
      17'd8267: data = 8'hfc;
      17'd8268: data = 8'hfc;
      17'd8269: data = 8'hf9;
      17'd8270: data = 8'hfe;
      17'd8271: data = 8'hfc;
      17'd8272: data = 8'hfd;
      17'd8273: data = 8'hfd;
      17'd8274: data = 8'hfd;
      17'd8275: data = 8'hfc;
      17'd8276: data = 8'hfc;
      17'd8277: data = 8'hfd;
      17'd8278: data = 8'hfc;
      17'd8279: data = 8'hfc;
      17'd8280: data = 8'hfe;
      17'd8281: data = 8'hfd;
      17'd8282: data = 8'hfc;
      17'd8283: data = 8'h00;
      17'd8284: data = 8'hfe;
      17'd8285: data = 8'hfd;
      17'd8286: data = 8'hfd;
      17'd8287: data = 8'hfc;
      17'd8288: data = 8'hfa;
      17'd8289: data = 8'hfd;
      17'd8290: data = 8'hfe;
      17'd8291: data = 8'hfe;
      17'd8292: data = 8'h01;
      17'd8293: data = 8'h02;
      17'd8294: data = 8'h00;
      17'd8295: data = 8'hfd;
      17'd8296: data = 8'hfe;
      17'd8297: data = 8'hfd;
      17'd8298: data = 8'h00;
      17'd8299: data = 8'hfd;
      17'd8300: data = 8'hfd;
      17'd8301: data = 8'h00;
      17'd8302: data = 8'h00;
      17'd8303: data = 8'h01;
      17'd8304: data = 8'h02;
      17'd8305: data = 8'h01;
      17'd8306: data = 8'h02;
      17'd8307: data = 8'h01;
      17'd8308: data = 8'hfe;
      17'd8309: data = 8'hfe;
      17'd8310: data = 8'h01;
      17'd8311: data = 8'h05;
      17'd8312: data = 8'h02;
      17'd8313: data = 8'h02;
      17'd8314: data = 8'h01;
      17'd8315: data = 8'h01;
      17'd8316: data = 8'h00;
      17'd8317: data = 8'h01;
      17'd8318: data = 8'h01;
      17'd8319: data = 8'hfe;
      17'd8320: data = 8'hfd;
      17'd8321: data = 8'h01;
      17'd8322: data = 8'h02;
      17'd8323: data = 8'h00;
      17'd8324: data = 8'hfe;
      17'd8325: data = 8'h00;
      17'd8326: data = 8'hfe;
      17'd8327: data = 8'hfd;
      17'd8328: data = 8'hfe;
      17'd8329: data = 8'hfc;
      17'd8330: data = 8'hfa;
      17'd8331: data = 8'hfe;
      17'd8332: data = 8'hfe;
      17'd8333: data = 8'hfe;
      17'd8334: data = 8'h00;
      17'd8335: data = 8'hfc;
      17'd8336: data = 8'hf9;
      17'd8337: data = 8'hfd;
      17'd8338: data = 8'h01;
      17'd8339: data = 8'hfa;
      17'd8340: data = 8'hf9;
      17'd8341: data = 8'h00;
      17'd8342: data = 8'h01;
      17'd8343: data = 8'hfe;
      17'd8344: data = 8'hfe;
      17'd8345: data = 8'h02;
      17'd8346: data = 8'h00;
      17'd8347: data = 8'hfa;
      17'd8348: data = 8'hfc;
      17'd8349: data = 8'h00;
      17'd8350: data = 8'hf9;
      17'd8351: data = 8'hfc;
      17'd8352: data = 8'h04;
      17'd8353: data = 8'h00;
      17'd8354: data = 8'hfc;
      17'd8355: data = 8'h01;
      17'd8356: data = 8'hfe;
      17'd8357: data = 8'hfc;
      17'd8358: data = 8'hfc;
      17'd8359: data = 8'h01;
      17'd8360: data = 8'h05;
      17'd8361: data = 8'h02;
      17'd8362: data = 8'h05;
      17'd8363: data = 8'hf6;
      17'd8364: data = 8'hf4;
      17'd8365: data = 8'hfa;
      17'd8366: data = 8'hfc;
      17'd8367: data = 8'hfc;
      17'd8368: data = 8'h01;
      17'd8369: data = 8'h05;
      17'd8370: data = 8'h05;
      17'd8371: data = 8'h05;
      17'd8372: data = 8'h0e;
      17'd8373: data = 8'h0a;
      17'd8374: data = 8'hfd;
      17'd8375: data = 8'hfc;
      17'd8376: data = 8'hf9;
      17'd8377: data = 8'hfa;
      17'd8378: data = 8'hfc;
      17'd8379: data = 8'hfd;
      17'd8380: data = 8'h00;
      17'd8381: data = 8'h11;
      17'd8382: data = 8'h0e;
      17'd8383: data = 8'h0c;
      17'd8384: data = 8'h0c;
      17'd8385: data = 8'hfe;
      17'd8386: data = 8'hf4;
      17'd8387: data = 8'hef;
      17'd8388: data = 8'hf4;
      17'd8389: data = 8'hf9;
      17'd8390: data = 8'h04;
      17'd8391: data = 8'h0e;
      17'd8392: data = 8'h0d;
      17'd8393: data = 8'h09;
      17'd8394: data = 8'h0c;
      17'd8395: data = 8'h04;
      17'd8396: data = 8'hfd;
      17'd8397: data = 8'hf5;
      17'd8398: data = 8'hf9;
      17'd8399: data = 8'hf4;
      17'd8400: data = 8'hfa;
      17'd8401: data = 8'h0d;
      17'd8402: data = 8'h15;
      17'd8403: data = 8'h0e;
      17'd8404: data = 8'h04;
      17'd8405: data = 8'hfe;
      17'd8406: data = 8'hf2;
      17'd8407: data = 8'hf1;
      17'd8408: data = 8'hf5;
      17'd8409: data = 8'hfd;
      17'd8410: data = 8'h09;
      17'd8411: data = 8'h0d;
      17'd8412: data = 8'h06;
      17'd8413: data = 8'h09;
      17'd8414: data = 8'h09;
      17'd8415: data = 8'hf9;
      17'd8416: data = 8'he0;
      17'd8417: data = 8'he5;
      17'd8418: data = 8'hfa;
      17'd8419: data = 8'h0a;
      17'd8420: data = 8'h16;
      17'd8421: data = 8'h19;
      17'd8422: data = 8'h09;
      17'd8423: data = 8'hf9;
      17'd8424: data = 8'hed;
      17'd8425: data = 8'he4;
      17'd8426: data = 8'he7;
      17'd8427: data = 8'hf9;
      17'd8428: data = 8'h09;
      17'd8429: data = 8'h12;
      17'd8430: data = 8'h19;
      17'd8431: data = 8'h19;
      17'd8432: data = 8'h11;
      17'd8433: data = 8'hfc;
      17'd8434: data = 8'hec;
      17'd8435: data = 8'he4;
      17'd8436: data = 8'he5;
      17'd8437: data = 8'hef;
      17'd8438: data = 8'h06;
      17'd8439: data = 8'h1a;
      17'd8440: data = 8'h1b;
      17'd8441: data = 8'h12;
      17'd8442: data = 8'h05;
      17'd8443: data = 8'hfc;
      17'd8444: data = 8'hf2;
      17'd8445: data = 8'hf2;
      17'd8446: data = 8'hf4;
      17'd8447: data = 8'hfa;
      17'd8448: data = 8'h0a;
      17'd8449: data = 8'h15;
      17'd8450: data = 8'h0e;
      17'd8451: data = 8'h06;
      17'd8452: data = 8'hfa;
      17'd8453: data = 8'hf5;
      17'd8454: data = 8'hf2;
      17'd8455: data = 8'hf1;
      17'd8456: data = 8'hf5;
      17'd8457: data = 8'hfa;
      17'd8458: data = 8'h0a;
      17'd8459: data = 8'h06;
      17'd8460: data = 8'h02;
      17'd8461: data = 8'h09;
      17'd8462: data = 8'hfd;
      17'd8463: data = 8'hed;
      17'd8464: data = 8'hed;
      17'd8465: data = 8'hf6;
      17'd8466: data = 8'h00;
      17'd8467: data = 8'h02;
      17'd8468: data = 8'h04;
      17'd8469: data = 8'h02;
      17'd8470: data = 8'h01;
      17'd8471: data = 8'hfc;
      17'd8472: data = 8'hf5;
      17'd8473: data = 8'hf1;
      17'd8474: data = 8'hf6;
      17'd8475: data = 8'hfa;
      17'd8476: data = 8'h01;
      17'd8477: data = 8'h06;
      17'd8478: data = 8'h0c;
      17'd8479: data = 8'h06;
      17'd8480: data = 8'hfc;
      17'd8481: data = 8'hfc;
      17'd8482: data = 8'hf6;
      17'd8483: data = 8'hef;
      17'd8484: data = 8'hf2;
      17'd8485: data = 8'hfc;
      17'd8486: data = 8'hfe;
      17'd8487: data = 8'h09;
      17'd8488: data = 8'h0e;
      17'd8489: data = 8'h06;
      17'd8490: data = 8'h04;
      17'd8491: data = 8'hfe;
      17'd8492: data = 8'hf5;
      17'd8493: data = 8'hf2;
      17'd8494: data = 8'hf5;
      17'd8495: data = 8'hfa;
      17'd8496: data = 8'h04;
      17'd8497: data = 8'h05;
      17'd8498: data = 8'h02;
      17'd8499: data = 8'hfe;
      17'd8500: data = 8'h01;
      17'd8501: data = 8'hfd;
      17'd8502: data = 8'hfa;
      17'd8503: data = 8'hfa;
      17'd8504: data = 8'hf6;
      17'd8505: data = 8'hfd;
      17'd8506: data = 8'h01;
      17'd8507: data = 8'h05;
      17'd8508: data = 8'h01;
      17'd8509: data = 8'hfc;
      17'd8510: data = 8'hf5;
      17'd8511: data = 8'hf6;
      17'd8512: data = 8'hf4;
      17'd8513: data = 8'hfd;
      17'd8514: data = 8'h0a;
      17'd8515: data = 8'h01;
      17'd8516: data = 8'hf6;
      17'd8517: data = 8'hed;
      17'd8518: data = 8'he9;
      17'd8519: data = 8'hf4;
      17'd8520: data = 8'hfd;
      17'd8521: data = 8'h01;
      17'd8522: data = 8'h01;
      17'd8523: data = 8'h00;
      17'd8524: data = 8'h01;
      17'd8525: data = 8'hf9;
      17'd8526: data = 8'hec;
      17'd8527: data = 8'heb;
      17'd8528: data = 8'hf4;
      17'd8529: data = 8'hfa;
      17'd8530: data = 8'hf9;
      17'd8531: data = 8'hfe;
      17'd8532: data = 8'h02;
      17'd8533: data = 8'h05;
      17'd8534: data = 8'h05;
      17'd8535: data = 8'hf2;
      17'd8536: data = 8'he7;
      17'd8537: data = 8'hef;
      17'd8538: data = 8'hfe;
      17'd8539: data = 8'h04;
      17'd8540: data = 8'h0a;
      17'd8541: data = 8'h13;
      17'd8542: data = 8'h11;
      17'd8543: data = 8'hfd;
      17'd8544: data = 8'hef;
      17'd8545: data = 8'hfc;
      17'd8546: data = 8'hf6;
      17'd8547: data = 8'hf9;
      17'd8548: data = 8'h0e;
      17'd8549: data = 8'h16;
      17'd8550: data = 8'h06;
      17'd8551: data = 8'h11;
      17'd8552: data = 8'h09;
      17'd8553: data = 8'h00;
      17'd8554: data = 8'h02;
      17'd8555: data = 8'hf9;
      17'd8556: data = 8'h01;
      17'd8557: data = 8'h09;
      17'd8558: data = 8'h0c;
      17'd8559: data = 8'h04;
      17'd8560: data = 8'h00;
      17'd8561: data = 8'h0e;
      17'd8562: data = 8'h0d;
      17'd8563: data = 8'h11;
      17'd8564: data = 8'h13;
      17'd8565: data = 8'hfc;
      17'd8566: data = 8'hf5;
      17'd8567: data = 8'hfd;
      17'd8568: data = 8'h02;
      17'd8569: data = 8'h15;
      17'd8570: data = 8'h1b;
      17'd8571: data = 8'h01;
      17'd8572: data = 8'hf5;
      17'd8573: data = 8'hf5;
      17'd8574: data = 8'hfc;
      17'd8575: data = 8'h16;
      17'd8576: data = 8'h13;
      17'd8577: data = 8'h0e;
      17'd8578: data = 8'h0a;
      17'd8579: data = 8'hf6;
      17'd8580: data = 8'hf1;
      17'd8581: data = 8'hec;
      17'd8582: data = 8'hec;
      17'd8583: data = 8'hf5;
      17'd8584: data = 8'h09;
      17'd8585: data = 8'h0a;
      17'd8586: data = 8'h11;
      17'd8587: data = 8'h0e;
      17'd8588: data = 8'h01;
      17'd8589: data = 8'hf6;
      17'd8590: data = 8'hf1;
      17'd8591: data = 8'hef;
      17'd8592: data = 8'he7;
      17'd8593: data = 8'hef;
      17'd8594: data = 8'h00;
      17'd8595: data = 8'h02;
      17'd8596: data = 8'hfd;
      17'd8597: data = 8'h0c;
      17'd8598: data = 8'h15;
      17'd8599: data = 8'hf5;
      17'd8600: data = 8'hef;
      17'd8601: data = 8'hef;
      17'd8602: data = 8'he5;
      17'd8603: data = 8'hf9;
      17'd8604: data = 8'h0a;
      17'd8605: data = 8'h09;
      17'd8606: data = 8'hf4;
      17'd8607: data = 8'hf2;
      17'd8608: data = 8'h00;
      17'd8609: data = 8'hf2;
      17'd8610: data = 8'hf4;
      17'd8611: data = 8'h16;
      17'd8612: data = 8'h0a;
      17'd8613: data = 8'he9;
      17'd8614: data = 8'he7;
      17'd8615: data = 8'hfc;
      17'd8616: data = 8'hfe;
      17'd8617: data = 8'hef;
      17'd8618: data = 8'hf5;
      17'd8619: data = 8'hfe;
      17'd8620: data = 8'hfd;
      17'd8621: data = 8'h04;
      17'd8622: data = 8'h02;
      17'd8623: data = 8'hfd;
      17'd8624: data = 8'h00;
      17'd8625: data = 8'hfc;
      17'd8626: data = 8'hf6;
      17'd8627: data = 8'hf5;
      17'd8628: data = 8'hfa;
      17'd8629: data = 8'hfd;
      17'd8630: data = 8'hfd;
      17'd8631: data = 8'hfd;
      17'd8632: data = 8'h05;
      17'd8633: data = 8'h0c;
      17'd8634: data = 8'h04;
      17'd8635: data = 8'h01;
      17'd8636: data = 8'h04;
      17'd8637: data = 8'hfe;
      17'd8638: data = 8'hf5;
      17'd8639: data = 8'hfc;
      17'd8640: data = 8'h0a;
      17'd8641: data = 8'h0a;
      17'd8642: data = 8'h04;
      17'd8643: data = 8'h09;
      17'd8644: data = 8'h0e;
      17'd8645: data = 8'h0c;
      17'd8646: data = 8'h0c;
      17'd8647: data = 8'h0c;
      17'd8648: data = 8'h04;
      17'd8649: data = 8'h01;
      17'd8650: data = 8'h04;
      17'd8651: data = 8'h06;
      17'd8652: data = 8'h0c;
      17'd8653: data = 8'h12;
      17'd8654: data = 8'h0c;
      17'd8655: data = 8'h09;
      17'd8656: data = 8'h0e;
      17'd8657: data = 8'h0a;
      17'd8658: data = 8'h06;
      17'd8659: data = 8'h0d;
      17'd8660: data = 8'h01;
      17'd8661: data = 8'hfa;
      17'd8662: data = 8'h00;
      17'd8663: data = 8'h02;
      17'd8664: data = 8'h05;
      17'd8665: data = 8'h04;
      17'd8666: data = 8'h06;
      17'd8667: data = 8'h01;
      17'd8668: data = 8'hfd;
      17'd8669: data = 8'hfe;
      17'd8670: data = 8'hfa;
      17'd8671: data = 8'hf6;
      17'd8672: data = 8'hf6;
      17'd8673: data = 8'hf2;
      17'd8674: data = 8'hfa;
      17'd8675: data = 8'h02;
      17'd8676: data = 8'hfc;
      17'd8677: data = 8'hfd;
      17'd8678: data = 8'hfe;
      17'd8679: data = 8'hfd;
      17'd8680: data = 8'hf9;
      17'd8681: data = 8'hf5;
      17'd8682: data = 8'hf6;
      17'd8683: data = 8'hf5;
      17'd8684: data = 8'hf4;
      17'd8685: data = 8'hfa;
      17'd8686: data = 8'hf6;
      17'd8687: data = 8'hfa;
      17'd8688: data = 8'hfe;
      17'd8689: data = 8'hfc;
      17'd8690: data = 8'hf9;
      17'd8691: data = 8'hfa;
      17'd8692: data = 8'h01;
      17'd8693: data = 8'h00;
      17'd8694: data = 8'hfa;
      17'd8695: data = 8'hf9;
      17'd8696: data = 8'hf5;
      17'd8697: data = 8'hf9;
      17'd8698: data = 8'h04;
      17'd8699: data = 8'h09;
      17'd8700: data = 8'h05;
      17'd8701: data = 8'h09;
      17'd8702: data = 8'h06;
      17'd8703: data = 8'hfc;
      17'd8704: data = 8'hf6;
      17'd8705: data = 8'h09;
      17'd8706: data = 8'h19;
      17'd8707: data = 8'h0e;
      17'd8708: data = 8'h05;
      17'd8709: data = 8'h0a;
      17'd8710: data = 8'h0a;
      17'd8711: data = 8'h0a;
      17'd8712: data = 8'h11;
      17'd8713: data = 8'h13;
      17'd8714: data = 8'h15;
      17'd8715: data = 8'h1f;
      17'd8716: data = 8'h16;
      17'd8717: data = 8'h06;
      17'd8718: data = 8'h05;
      17'd8719: data = 8'h0d;
      17'd8720: data = 8'h11;
      17'd8721: data = 8'h11;
      17'd8722: data = 8'h1b;
      17'd8723: data = 8'h24;
      17'd8724: data = 8'h1a;
      17'd8725: data = 8'h11;
      17'd8726: data = 8'h0c;
      17'd8727: data = 8'h09;
      17'd8728: data = 8'h0e;
      17'd8729: data = 8'h12;
      17'd8730: data = 8'h0c;
      17'd8731: data = 8'h0d;
      17'd8732: data = 8'h0a;
      17'd8733: data = 8'h02;
      17'd8734: data = 8'h0a;
      17'd8735: data = 8'h15;
      17'd8736: data = 8'h0e;
      17'd8737: data = 8'h0a;
      17'd8738: data = 8'h01;
      17'd8739: data = 8'hf4;
      17'd8740: data = 8'hfd;
      17'd8741: data = 8'h04;
      17'd8742: data = 8'h02;
      17'd8743: data = 8'h01;
      17'd8744: data = 8'h00;
      17'd8745: data = 8'hf9;
      17'd8746: data = 8'hf2;
      17'd8747: data = 8'hed;
      17'd8748: data = 8'hf9;
      17'd8749: data = 8'hfd;
      17'd8750: data = 8'hed;
      17'd8751: data = 8'hec;
      17'd8752: data = 8'hef;
      17'd8753: data = 8'hed;
      17'd8754: data = 8'he7;
      17'd8755: data = 8'he4;
      17'd8756: data = 8'he3;
      17'd8757: data = 8'he0;
      17'd8758: data = 8'he7;
      17'd8759: data = 8'hef;
      17'd8760: data = 8'hdb;
      17'd8761: data = 8'hdb;
      17'd8762: data = 8'hd3;
      17'd8763: data = 8'hd1;
      17'd8764: data = 8'hda;
      17'd8765: data = 8'hde;
      17'd8766: data = 8'heb;
      17'd8767: data = 8'he2;
      17'd8768: data = 8'hcd;
      17'd8769: data = 8'hd5;
      17'd8770: data = 8'hef;
      17'd8771: data = 8'he2;
      17'd8772: data = 8'hda;
      17'd8773: data = 8'he5;
      17'd8774: data = 8'hdb;
      17'd8775: data = 8'hd3;
      17'd8776: data = 8'hf2;
      17'd8777: data = 8'h01;
      17'd8778: data = 8'hf2;
      17'd8779: data = 8'hdb;
      17'd8780: data = 8'hdc;
      17'd8781: data = 8'hf2;
      17'd8782: data = 8'hfa;
      17'd8783: data = 8'h00;
      17'd8784: data = 8'hf6;
      17'd8785: data = 8'hf5;
      17'd8786: data = 8'hf2;
      17'd8787: data = 8'hfa;
      17'd8788: data = 8'hfd;
      17'd8789: data = 8'h05;
      17'd8790: data = 8'h11;
      17'd8791: data = 8'h09;
      17'd8792: data = 8'hfe;
      17'd8793: data = 8'hfe;
      17'd8794: data = 8'h06;
      17'd8795: data = 8'h05;
      17'd8796: data = 8'h09;
      17'd8797: data = 8'hfa;
      17'd8798: data = 8'h01;
      17'd8799: data = 8'h0a;
      17'd8800: data = 8'h0c;
      17'd8801: data = 8'h15;
      17'd8802: data = 8'h16;
      17'd8803: data = 8'h13;
      17'd8804: data = 8'h00;
      17'd8805: data = 8'hfa;
      17'd8806: data = 8'h0a;
      17'd8807: data = 8'h11;
      17'd8808: data = 8'h0e;
      17'd8809: data = 8'h0e;
      17'd8810: data = 8'h16;
      17'd8811: data = 8'h0a;
      17'd8812: data = 8'hf6;
      17'd8813: data = 8'hfe;
      17'd8814: data = 8'h05;
      17'd8815: data = 8'h01;
      17'd8816: data = 8'h09;
      17'd8817: data = 8'h12;
      17'd8818: data = 8'h0c;
      17'd8819: data = 8'h0a;
      17'd8820: data = 8'hfd;
      17'd8821: data = 8'hed;
      17'd8822: data = 8'hef;
      17'd8823: data = 8'h01;
      17'd8824: data = 8'h0e;
      17'd8825: data = 8'h0e;
      17'd8826: data = 8'h0d;
      17'd8827: data = 8'hf4;
      17'd8828: data = 8'hed;
      17'd8829: data = 8'hf2;
      17'd8830: data = 8'hf5;
      17'd8831: data = 8'h09;
      17'd8832: data = 8'h13;
      17'd8833: data = 8'h0c;
      17'd8834: data = 8'hfc;
      17'd8835: data = 8'hf6;
      17'd8836: data = 8'hfd;
      17'd8837: data = 8'h04;
      17'd8838: data = 8'h06;
      17'd8839: data = 8'h01;
      17'd8840: data = 8'hfe;
      17'd8841: data = 8'h01;
      17'd8842: data = 8'h00;
      17'd8843: data = 8'hfe;
      17'd8844: data = 8'h09;
      17'd8845: data = 8'h0c;
      17'd8846: data = 8'h05;
      17'd8847: data = 8'h05;
      17'd8848: data = 8'h05;
      17'd8849: data = 8'h0a;
      17'd8850: data = 8'h11;
      17'd8851: data = 8'h11;
      17'd8852: data = 8'h09;
      17'd8853: data = 8'h09;
      17'd8854: data = 8'h13;
      17'd8855: data = 8'h12;
      17'd8856: data = 8'h04;
      17'd8857: data = 8'h06;
      17'd8858: data = 8'h11;
      17'd8859: data = 8'h0e;
      17'd8860: data = 8'h12;
      17'd8861: data = 8'h15;
      17'd8862: data = 8'h16;
      17'd8863: data = 8'h0e;
      17'd8864: data = 8'h06;
      17'd8865: data = 8'h09;
      17'd8866: data = 8'h11;
      17'd8867: data = 8'h16;
      17'd8868: data = 8'h13;
      17'd8869: data = 8'h06;
      17'd8870: data = 8'h02;
      17'd8871: data = 8'h05;
      17'd8872: data = 8'h0a;
      17'd8873: data = 8'h09;
      17'd8874: data = 8'h02;
      17'd8875: data = 8'h01;
      17'd8876: data = 8'h02;
      17'd8877: data = 8'h01;
      17'd8878: data = 8'hfd;
      17'd8879: data = 8'h01;
      17'd8880: data = 8'h04;
      17'd8881: data = 8'hfd;
      17'd8882: data = 8'hf6;
      17'd8883: data = 8'hfc;
      17'd8884: data = 8'hfe;
      17'd8885: data = 8'hfd;
      17'd8886: data = 8'hfa;
      17'd8887: data = 8'hf9;
      17'd8888: data = 8'hf9;
      17'd8889: data = 8'hfa;
      17'd8890: data = 8'hfa;
      17'd8891: data = 8'hfc;
      17'd8892: data = 8'hfc;
      17'd8893: data = 8'hfd;
      17'd8894: data = 8'hfd;
      17'd8895: data = 8'hf6;
      17'd8896: data = 8'hf5;
      17'd8897: data = 8'hfe;
      17'd8898: data = 8'h02;
      17'd8899: data = 8'hfc;
      17'd8900: data = 8'hfa;
      17'd8901: data = 8'h04;
      17'd8902: data = 8'h05;
      17'd8903: data = 8'h04;
      17'd8904: data = 8'h02;
      17'd8905: data = 8'h00;
      17'd8906: data = 8'h04;
      17'd8907: data = 8'h04;
      17'd8908: data = 8'h06;
      17'd8909: data = 8'h0c;
      17'd8910: data = 8'h09;
      17'd8911: data = 8'h0a;
      17'd8912: data = 8'h09;
      17'd8913: data = 8'h05;
      17'd8914: data = 8'h0d;
      17'd8915: data = 8'h11;
      17'd8916: data = 8'h0d;
      17'd8917: data = 8'h0a;
      17'd8918: data = 8'h0c;
      17'd8919: data = 8'h12;
      17'd8920: data = 8'h12;
      17'd8921: data = 8'h0a;
      17'd8922: data = 8'h02;
      17'd8923: data = 8'h09;
      17'd8924: data = 8'h12;
      17'd8925: data = 8'h12;
      17'd8926: data = 8'h0c;
      17'd8927: data = 8'h0c;
      17'd8928: data = 8'h0d;
      17'd8929: data = 8'h06;
      17'd8930: data = 8'h02;
      17'd8931: data = 8'h04;
      17'd8932: data = 8'h15;
      17'd8933: data = 8'h15;
      17'd8934: data = 8'h0d;
      17'd8935: data = 8'h13;
      17'd8936: data = 8'h05;
      17'd8937: data = 8'h00;
      17'd8938: data = 8'h01;
      17'd8939: data = 8'h02;
      17'd8940: data = 8'h05;
      17'd8941: data = 8'h0d;
      17'd8942: data = 8'h11;
      17'd8943: data = 8'h06;
      17'd8944: data = 8'h04;
      17'd8945: data = 8'h04;
      17'd8946: data = 8'hfc;
      17'd8947: data = 8'hf9;
      17'd8948: data = 8'h01;
      17'd8949: data = 8'h0d;
      17'd8950: data = 8'h0c;
      17'd8951: data = 8'hfa;
      17'd8952: data = 8'hf4;
      17'd8953: data = 8'hf6;
      17'd8954: data = 8'hf9;
      17'd8955: data = 8'hf9;
      17'd8956: data = 8'hf6;
      17'd8957: data = 8'hf5;
      17'd8958: data = 8'hf5;
      17'd8959: data = 8'hf9;
      17'd8960: data = 8'hf5;
      17'd8961: data = 8'hf1;
      17'd8962: data = 8'heb;
      17'd8963: data = 8'hef;
      17'd8964: data = 8'hf2;
      17'd8965: data = 8'heb;
      17'd8966: data = 8'he9;
      17'd8967: data = 8'heb;
      17'd8968: data = 8'he9;
      17'd8969: data = 8'hde;
      17'd8970: data = 8'hde;
      17'd8971: data = 8'he2;
      17'd8972: data = 8'hd5;
      17'd8973: data = 8'hdb;
      17'd8974: data = 8'he4;
      17'd8975: data = 8'he7;
      17'd8976: data = 8'he7;
      17'd8977: data = 8'hda;
      17'd8978: data = 8'hd5;
      17'd8979: data = 8'hd2;
      17'd8980: data = 8'hda;
      17'd8981: data = 8'hd5;
      17'd8982: data = 8'hd2;
      17'd8983: data = 8'hdb;
      17'd8984: data = 8'hde;
      17'd8985: data = 8'hda;
      17'd8986: data = 8'hd6;
      17'd8987: data = 8'hd3;
      17'd8988: data = 8'hd6;
      17'd8989: data = 8'hde;
      17'd8990: data = 8'he5;
      17'd8991: data = 8'he7;
      17'd8992: data = 8'he3;
      17'd8993: data = 8'he2;
      17'd8994: data = 8'hd6;
      17'd8995: data = 8'hd6;
      17'd8996: data = 8'he7;
      17'd8997: data = 8'hfd;
      17'd8998: data = 8'hfd;
      17'd8999: data = 8'hf6;
      17'd9000: data = 8'hec;
      17'd9001: data = 8'he3;
      17'd9002: data = 8'he7;
      17'd9003: data = 8'hf2;
      17'd9004: data = 8'hfe;
      17'd9005: data = 8'h04;
      17'd9006: data = 8'h0e;
      17'd9007: data = 8'h06;
      17'd9008: data = 8'h04;
      17'd9009: data = 8'hfe;
      17'd9010: data = 8'h0a;
      17'd9011: data = 8'h0c;
      17'd9012: data = 8'h06;
      17'd9013: data = 8'h15;
      17'd9014: data = 8'h15;
      17'd9015: data = 8'h15;
      17'd9016: data = 8'h12;
      17'd9017: data = 8'h0d;
      17'd9018: data = 8'h05;
      17'd9019: data = 8'h0e;
      17'd9020: data = 8'h13;
      17'd9021: data = 8'h12;
      17'd9022: data = 8'h19;
      17'd9023: data = 8'h22;
      17'd9024: data = 8'h1f;
      17'd9025: data = 8'h0e;
      17'd9026: data = 8'h11;
      17'd9027: data = 8'h12;
      17'd9028: data = 8'h0d;
      17'd9029: data = 8'h0c;
      17'd9030: data = 8'h0e;
      17'd9031: data = 8'h1c;
      17'd9032: data = 8'h24;
      17'd9033: data = 8'h11;
      17'd9034: data = 8'h01;
      17'd9035: data = 8'h02;
      17'd9036: data = 8'h09;
      17'd9037: data = 8'h0c;
      17'd9038: data = 8'h16;
      17'd9039: data = 8'h1a;
      17'd9040: data = 8'h0c;
      17'd9041: data = 8'h0c;
      17'd9042: data = 8'h01;
      17'd9043: data = 8'hf2;
      17'd9044: data = 8'hf9;
      17'd9045: data = 8'h06;
      17'd9046: data = 8'h0a;
      17'd9047: data = 8'h0a;
      17'd9048: data = 8'h15;
      17'd9049: data = 8'h05;
      17'd9050: data = 8'hec;
      17'd9051: data = 8'he4;
      17'd9052: data = 8'heb;
      17'd9053: data = 8'hfe;
      17'd9054: data = 8'h16;
      17'd9055: data = 8'h1e;
      17'd9056: data = 8'h15;
      17'd9057: data = 8'h01;
      17'd9058: data = 8'hef;
      17'd9059: data = 8'he7;
      17'd9060: data = 8'hf1;
      17'd9061: data = 8'h01;
      17'd9062: data = 8'h11;
      17'd9063: data = 8'h1c;
      17'd9064: data = 8'h11;
      17'd9065: data = 8'hfc;
      17'd9066: data = 8'hf6;
      17'd9067: data = 8'hf6;
      17'd9068: data = 8'hf9;
      17'd9069: data = 8'h04;
      17'd9070: data = 8'h19;
      17'd9071: data = 8'h1e;
      17'd9072: data = 8'h16;
      17'd9073: data = 8'h04;
      17'd9074: data = 8'hf5;
      17'd9075: data = 8'hfd;
      17'd9076: data = 8'h04;
      17'd9077: data = 8'h11;
      17'd9078: data = 8'h1c;
      17'd9079: data = 8'h1b;
      17'd9080: data = 8'h11;
      17'd9081: data = 8'h04;
      17'd9082: data = 8'hfd;
      17'd9083: data = 8'h05;
      17'd9084: data = 8'h19;
      17'd9085: data = 8'h1c;
      17'd9086: data = 8'h16;
      17'd9087: data = 8'h0d;
      17'd9088: data = 8'h06;
      17'd9089: data = 8'h05;
      17'd9090: data = 8'h05;
      17'd9091: data = 8'h09;
      17'd9092: data = 8'h12;
      17'd9093: data = 8'h0e;
      17'd9094: data = 8'h04;
      17'd9095: data = 8'hfe;
      17'd9096: data = 8'hf9;
      17'd9097: data = 8'hfe;
      17'd9098: data = 8'h05;
      17'd9099: data = 8'h05;
      17'd9100: data = 8'h04;
      17'd9101: data = 8'h04;
      17'd9102: data = 8'hfd;
      17'd9103: data = 8'hf6;
      17'd9104: data = 8'hf4;
      17'd9105: data = 8'hf5;
      17'd9106: data = 8'hfa;
      17'd9107: data = 8'hfd;
      17'd9108: data = 8'hf5;
      17'd9109: data = 8'hf1;
      17'd9110: data = 8'hf5;
      17'd9111: data = 8'hf4;
      17'd9112: data = 8'hf6;
      17'd9113: data = 8'hfc;
      17'd9114: data = 8'hfd;
      17'd9115: data = 8'hf6;
      17'd9116: data = 8'hf2;
      17'd9117: data = 8'hec;
      17'd9118: data = 8'hf2;
      17'd9119: data = 8'hfd;
      17'd9120: data = 8'hfd;
      17'd9121: data = 8'hfd;
      17'd9122: data = 8'hfc;
      17'd9123: data = 8'hf9;
      17'd9124: data = 8'hfa;
      17'd9125: data = 8'hfa;
      17'd9126: data = 8'hf6;
      17'd9127: data = 8'h04;
      17'd9128: data = 8'h09;
      17'd9129: data = 8'h01;
      17'd9130: data = 8'hfd;
      17'd9131: data = 8'hfc;
      17'd9132: data = 8'h01;
      17'd9133: data = 8'h04;
      17'd9134: data = 8'h02;
      17'd9135: data = 8'h05;
      17'd9136: data = 8'h0a;
      17'd9137: data = 8'h06;
      17'd9138: data = 8'h00;
      17'd9139: data = 8'h01;
      17'd9140: data = 8'h02;
      17'd9141: data = 8'h06;
      17'd9142: data = 8'h0e;
      17'd9143: data = 8'h0c;
      17'd9144: data = 8'h09;
      17'd9145: data = 8'h0c;
      17'd9146: data = 8'h09;
      17'd9147: data = 8'h02;
      17'd9148: data = 8'h02;
      17'd9149: data = 8'h00;
      17'd9150: data = 8'h0a;
      17'd9151: data = 8'h12;
      17'd9152: data = 8'h0c;
      17'd9153: data = 8'h0c;
      17'd9154: data = 8'h0a;
      17'd9155: data = 8'h04;
      17'd9156: data = 8'h04;
      17'd9157: data = 8'h06;
      17'd9158: data = 8'h09;
      17'd9159: data = 8'h0a;
      17'd9160: data = 8'h0a;
      17'd9161: data = 8'h04;
      17'd9162: data = 8'h09;
      17'd9163: data = 8'h09;
      17'd9164: data = 8'hfe;
      17'd9165: data = 8'hfe;
      17'd9166: data = 8'h02;
      17'd9167: data = 8'h09;
      17'd9168: data = 8'h05;
      17'd9169: data = 8'h02;
      17'd9170: data = 8'h04;
      17'd9171: data = 8'hfd;
      17'd9172: data = 8'h00;
      17'd9173: data = 8'h00;
      17'd9174: data = 8'hfd;
      17'd9175: data = 8'h00;
      17'd9176: data = 8'h00;
      17'd9177: data = 8'hfc;
      17'd9178: data = 8'hf4;
      17'd9179: data = 8'hf5;
      17'd9180: data = 8'hf6;
      17'd9181: data = 8'hfa;
      17'd9182: data = 8'hfd;
      17'd9183: data = 8'hf5;
      17'd9184: data = 8'hed;
      17'd9185: data = 8'hef;
      17'd9186: data = 8'heb;
      17'd9187: data = 8'heb;
      17'd9188: data = 8'hed;
      17'd9189: data = 8'hec;
      17'd9190: data = 8'he9;
      17'd9191: data = 8'he5;
      17'd9192: data = 8'he9;
      17'd9193: data = 8'he7;
      17'd9194: data = 8'he3;
      17'd9195: data = 8'hd6;
      17'd9196: data = 8'hd8;
      17'd9197: data = 8'he4;
      17'd9198: data = 8'hde;
      17'd9199: data = 8'hde;
      17'd9200: data = 8'hdb;
      17'd9201: data = 8'hd8;
      17'd9202: data = 8'hdc;
      17'd9203: data = 8'hda;
      17'd9204: data = 8'hd8;
      17'd9205: data = 8'hd8;
      17'd9206: data = 8'hdb;
      17'd9207: data = 8'hd8;
      17'd9208: data = 8'hd3;
      17'd9209: data = 8'hd3;
      17'd9210: data = 8'hdb;
      17'd9211: data = 8'hde;
      17'd9212: data = 8'hda;
      17'd9213: data = 8'hdb;
      17'd9214: data = 8'hd6;
      17'd9215: data = 8'he2;
      17'd9216: data = 8'he2;
      17'd9217: data = 8'hde;
      17'd9218: data = 8'he0;
      17'd9219: data = 8'he5;
      17'd9220: data = 8'he9;
      17'd9221: data = 8'hec;
      17'd9222: data = 8'hfa;
      17'd9223: data = 8'hf5;
      17'd9224: data = 8'hf1;
      17'd9225: data = 8'he5;
      17'd9226: data = 8'hef;
      17'd9227: data = 8'h0e;
      17'd9228: data = 8'h0e;
      17'd9229: data = 8'hfa;
      17'd9230: data = 8'hfa;
      17'd9231: data = 8'h0e;
      17'd9232: data = 8'h09;
      17'd9233: data = 8'hf6;
      17'd9234: data = 8'h0c;
      17'd9235: data = 8'h1b;
      17'd9236: data = 8'h12;
      17'd9237: data = 8'h16;
      17'd9238: data = 8'h1c;
      17'd9239: data = 8'h13;
      17'd9240: data = 8'h15;
      17'd9241: data = 8'h22;
      17'd9242: data = 8'h1f;
      17'd9243: data = 8'h1c;
      17'd9244: data = 8'h1e;
      17'd9245: data = 8'h1e;
      17'd9246: data = 8'h12;
      17'd9247: data = 8'h19;
      17'd9248: data = 8'h29;
      17'd9249: data = 8'h1f;
      17'd9250: data = 8'h23;
      17'd9251: data = 8'h27;
      17'd9252: data = 8'h1c;
      17'd9253: data = 8'h12;
      17'd9254: data = 8'h13;
      17'd9255: data = 8'h1f;
      17'd9256: data = 8'h1c;
      17'd9257: data = 8'h24;
      17'd9258: data = 8'h1c;
      17'd9259: data = 8'h11;
      17'd9260: data = 8'h12;
      17'd9261: data = 8'h16;
      17'd9262: data = 8'h0c;
      17'd9263: data = 8'h04;
      17'd9264: data = 8'h15;
      17'd9265: data = 8'h0d;
      17'd9266: data = 8'h06;
      17'd9267: data = 8'h12;
      17'd9268: data = 8'h12;
      17'd9269: data = 8'h0a;
      17'd9270: data = 8'hfd;
      17'd9271: data = 8'hfa;
      17'd9272: data = 8'h0a;
      17'd9273: data = 8'h02;
      17'd9274: data = 8'hfd;
      17'd9275: data = 8'h05;
      17'd9276: data = 8'h05;
      17'd9277: data = 8'h05;
      17'd9278: data = 8'hfd;
      17'd9279: data = 8'hf4;
      17'd9280: data = 8'heb;
      17'd9281: data = 8'hf1;
      17'd9282: data = 8'h06;
      17'd9283: data = 8'h11;
      17'd9284: data = 8'h12;
      17'd9285: data = 8'h0d;
      17'd9286: data = 8'hf5;
      17'd9287: data = 8'he2;
      17'd9288: data = 8'he3;
      17'd9289: data = 8'hfd;
      17'd9290: data = 8'h11;
      17'd9291: data = 8'h13;
      17'd9292: data = 8'h13;
      17'd9293: data = 8'hfc;
      17'd9294: data = 8'he7;
      17'd9295: data = 8'hed;
      17'd9296: data = 8'hf6;
      17'd9297: data = 8'h06;
      17'd9298: data = 8'h22;
      17'd9299: data = 8'h1c;
      17'd9300: data = 8'h06;
      17'd9301: data = 8'hfd;
      17'd9302: data = 8'hf4;
      17'd9303: data = 8'hf2;
      17'd9304: data = 8'hfe;
      17'd9305: data = 8'h13;
      17'd9306: data = 8'h23;
      17'd9307: data = 8'h1f;
      17'd9308: data = 8'h0d;
      17'd9309: data = 8'hf9;
      17'd9310: data = 8'hf1;
      17'd9311: data = 8'hfe;
      17'd9312: data = 8'h12;
      17'd9313: data = 8'h23;
      17'd9314: data = 8'h1e;
      17'd9315: data = 8'h0e;
      17'd9316: data = 8'h02;
      17'd9317: data = 8'hf6;
      17'd9318: data = 8'hfc;
      17'd9319: data = 8'h05;
      17'd9320: data = 8'h13;
      17'd9321: data = 8'h19;
      17'd9322: data = 8'h05;
      17'd9323: data = 8'hfc;
      17'd9324: data = 8'hfa;
      17'd9325: data = 8'hf9;
      17'd9326: data = 8'hfe;
      17'd9327: data = 8'h05;
      17'd9328: data = 8'h06;
      17'd9329: data = 8'h01;
      17'd9330: data = 8'hfd;
      17'd9331: data = 8'hf5;
      17'd9332: data = 8'hed;
      17'd9333: data = 8'hfa;
      17'd9334: data = 8'hfc;
      17'd9335: data = 8'hfc;
      17'd9336: data = 8'hfd;
      17'd9337: data = 8'hf6;
      17'd9338: data = 8'hf5;
      17'd9339: data = 8'hf5;
      17'd9340: data = 8'hed;
      17'd9341: data = 8'hf5;
      17'd9342: data = 8'hfc;
      17'd9343: data = 8'hf5;
      17'd9344: data = 8'hf5;
      17'd9345: data = 8'hf2;
      17'd9346: data = 8'hf2;
      17'd9347: data = 8'hfa;
      17'd9348: data = 8'hfd;
      17'd9349: data = 8'hfd;
      17'd9350: data = 8'hfc;
      17'd9351: data = 8'hf6;
      17'd9352: data = 8'hf1;
      17'd9353: data = 8'hf6;
      17'd9354: data = 8'hfc;
      17'd9355: data = 8'h00;
      17'd9356: data = 8'h01;
      17'd9357: data = 8'hfd;
      17'd9358: data = 8'hf6;
      17'd9359: data = 8'hfa;
      17'd9360: data = 8'h00;
      17'd9361: data = 8'h01;
      17'd9362: data = 8'h06;
      17'd9363: data = 8'h06;
      17'd9364: data = 8'h04;
      17'd9365: data = 8'hfe;
      17'd9366: data = 8'hf9;
      17'd9367: data = 8'h00;
      17'd9368: data = 8'h05;
      17'd9369: data = 8'h00;
      17'd9370: data = 8'h05;
      17'd9371: data = 8'h0a;
      17'd9372: data = 8'h06;
      17'd9373: data = 8'h04;
      17'd9374: data = 8'hfe;
      17'd9375: data = 8'hfa;
      17'd9376: data = 8'h04;
      17'd9377: data = 8'h11;
      17'd9378: data = 8'h0d;
      17'd9379: data = 8'h0c;
      17'd9380: data = 8'h0a;
      17'd9381: data = 8'hfc;
      17'd9382: data = 8'hf4;
      17'd9383: data = 8'h00;
      17'd9384: data = 8'h05;
      17'd9385: data = 8'h05;
      17'd9386: data = 8'h0e;
      17'd9387: data = 8'h15;
      17'd9388: data = 8'h06;
      17'd9389: data = 8'hfc;
      17'd9390: data = 8'h00;
      17'd9391: data = 8'hfd;
      17'd9392: data = 8'hfd;
      17'd9393: data = 8'h13;
      17'd9394: data = 8'h1b;
      17'd9395: data = 8'h06;
      17'd9396: data = 8'h00;
      17'd9397: data = 8'h01;
      17'd9398: data = 8'hf6;
      17'd9399: data = 8'hf5;
      17'd9400: data = 8'h01;
      17'd9401: data = 8'h06;
      17'd9402: data = 8'h0a;
      17'd9403: data = 8'h0a;
      17'd9404: data = 8'h00;
      17'd9405: data = 8'hf1;
      17'd9406: data = 8'hf2;
      17'd9407: data = 8'hfe;
      17'd9408: data = 8'h02;
      17'd9409: data = 8'h02;
      17'd9410: data = 8'hfd;
      17'd9411: data = 8'hf2;
      17'd9412: data = 8'hed;
      17'd9413: data = 8'hed;
      17'd9414: data = 8'hf1;
      17'd9415: data = 8'hf4;
      17'd9416: data = 8'hf5;
      17'd9417: data = 8'hf6;
      17'd9418: data = 8'hf4;
      17'd9419: data = 8'hef;
      17'd9420: data = 8'hec;
      17'd9421: data = 8'he3;
      17'd9422: data = 8'he3;
      17'd9423: data = 8'heb;
      17'd9424: data = 8'hec;
      17'd9425: data = 8'he9;
      17'd9426: data = 8'he2;
      17'd9427: data = 8'he4;
      17'd9428: data = 8'he5;
      17'd9429: data = 8'he0;
      17'd9430: data = 8'hdb;
      17'd9431: data = 8'hda;
      17'd9432: data = 8'he0;
      17'd9433: data = 8'he7;
      17'd9434: data = 8'he5;
      17'd9435: data = 8'hdc;
      17'd9436: data = 8'hd5;
      17'd9437: data = 8'hde;
      17'd9438: data = 8'hda;
      17'd9439: data = 8'hd2;
      17'd9440: data = 8'he3;
      17'd9441: data = 8'he4;
      17'd9442: data = 8'hdc;
      17'd9443: data = 8'hdb;
      17'd9444: data = 8'hdc;
      17'd9445: data = 8'hdb;
      17'd9446: data = 8'hda;
      17'd9447: data = 8'hdc;
      17'd9448: data = 8'he9;
      17'd9449: data = 8'hef;
      17'd9450: data = 8'hf4;
      17'd9451: data = 8'hf1;
      17'd9452: data = 8'he4;
      17'd9453: data = 8'he5;
      17'd9454: data = 8'hec;
      17'd9455: data = 8'h01;
      17'd9456: data = 8'hf6;
      17'd9457: data = 8'hf4;
      17'd9458: data = 8'h01;
      17'd9459: data = 8'hf9;
      17'd9460: data = 8'hfc;
      17'd9461: data = 8'h06;
      17'd9462: data = 8'h1b;
      17'd9463: data = 8'h04;
      17'd9464: data = 8'h00;
      17'd9465: data = 8'h1c;
      17'd9466: data = 8'h0d;
      17'd9467: data = 8'h12;
      17'd9468: data = 8'h1e;
      17'd9469: data = 8'h1b;
      17'd9470: data = 8'h16;
      17'd9471: data = 8'h16;
      17'd9472: data = 8'h1f;
      17'd9473: data = 8'h19;
      17'd9474: data = 8'h13;
      17'd9475: data = 8'h1f;
      17'd9476: data = 8'h23;
      17'd9477: data = 8'h1c;
      17'd9478: data = 8'h26;
      17'd9479: data = 8'h2c;
      17'd9480: data = 8'h1a;
      17'd9481: data = 8'h11;
      17'd9482: data = 8'h1f;
      17'd9483: data = 8'h1c;
      17'd9484: data = 8'h1b;
      17'd9485: data = 8'h29;
      17'd9486: data = 8'h29;
      17'd9487: data = 8'h1e;
      17'd9488: data = 8'h0d;
      17'd9489: data = 8'h06;
      17'd9490: data = 8'h15;
      17'd9491: data = 8'h16;
      17'd9492: data = 8'h26;
      17'd9493: data = 8'h1e;
      17'd9494: data = 8'h09;
      17'd9495: data = 8'h0c;
      17'd9496: data = 8'h12;
      17'd9497: data = 8'h0d;
      17'd9498: data = 8'h09;
      17'd9499: data = 8'h0e;
      17'd9500: data = 8'h0d;
      17'd9501: data = 8'h0e;
      17'd9502: data = 8'h15;
      17'd9503: data = 8'h09;
      17'd9504: data = 8'hf5;
      17'd9505: data = 8'hec;
      17'd9506: data = 8'hf9;
      17'd9507: data = 8'h04;
      17'd9508: data = 8'h0c;
      17'd9509: data = 8'h16;
      17'd9510: data = 8'h0a;
      17'd9511: data = 8'hf2;
      17'd9512: data = 8'hed;
      17'd9513: data = 8'hf1;
      17'd9514: data = 8'hf1;
      17'd9515: data = 8'h00;
      17'd9516: data = 8'h12;
      17'd9517: data = 8'h0e;
      17'd9518: data = 8'h02;
      17'd9519: data = 8'hf5;
      17'd9520: data = 8'he9;
      17'd9521: data = 8'he5;
      17'd9522: data = 8'hfd;
      17'd9523: data = 8'h05;
      17'd9524: data = 8'h04;
      17'd9525: data = 8'h0e;
      17'd9526: data = 8'h05;
      17'd9527: data = 8'hfc;
      17'd9528: data = 8'hf2;
      17'd9529: data = 8'hec;
      17'd9530: data = 8'hf6;
      17'd9531: data = 8'h15;
      17'd9532: data = 8'h24;
      17'd9533: data = 8'h15;
      17'd9534: data = 8'hfe;
      17'd9535: data = 8'hf1;
      17'd9536: data = 8'hed;
      17'd9537: data = 8'hf9;
      17'd9538: data = 8'h0d;
      17'd9539: data = 8'h1b;
      17'd9540: data = 8'h1c;
      17'd9541: data = 8'h11;
      17'd9542: data = 8'h01;
      17'd9543: data = 8'hfa;
      17'd9544: data = 8'hfa;
      17'd9545: data = 8'h06;
      17'd9546: data = 8'h15;
      17'd9547: data = 8'h1b;
      17'd9548: data = 8'h16;
      17'd9549: data = 8'h05;
      17'd9550: data = 8'hfc;
      17'd9551: data = 8'hf5;
      17'd9552: data = 8'hfc;
      17'd9553: data = 8'h0a;
      17'd9554: data = 8'h15;
      17'd9555: data = 8'h0d;
      17'd9556: data = 8'h05;
      17'd9557: data = 8'h06;
      17'd9558: data = 8'hfa;
      17'd9559: data = 8'hf1;
      17'd9560: data = 8'hf5;
      17'd9561: data = 8'hfe;
      17'd9562: data = 8'h06;
      17'd9563: data = 8'h0a;
      17'd9564: data = 8'hfc;
      17'd9565: data = 8'hed;
      17'd9566: data = 8'hed;
      17'd9567: data = 8'hf4;
      17'd9568: data = 8'hfc;
      17'd9569: data = 8'hfc;
      17'd9570: data = 8'hf9;
      17'd9571: data = 8'hfc;
      17'd9572: data = 8'hf9;
      17'd9573: data = 8'hef;
      17'd9574: data = 8'hf4;
      17'd9575: data = 8'hfa;
      17'd9576: data = 8'hf5;
      17'd9577: data = 8'hf2;
      17'd9578: data = 8'hf5;
      17'd9579: data = 8'hf6;
      17'd9580: data = 8'hf4;
      17'd9581: data = 8'hf2;
      17'd9582: data = 8'hf5;
      17'd9583: data = 8'hfa;
      17'd9584: data = 8'hfc;
      17'd9585: data = 8'hf6;
      17'd9586: data = 8'hf5;
      17'd9587: data = 8'hfd;
      17'd9588: data = 8'h01;
      17'd9589: data = 8'h04;
      17'd9590: data = 8'hfd;
      17'd9591: data = 8'hfa;
      17'd9592: data = 8'hfc;
      17'd9593: data = 8'hfe;
      17'd9594: data = 8'h00;
      17'd9595: data = 8'hfe;
      17'd9596: data = 8'h01;
      17'd9597: data = 8'h02;
      17'd9598: data = 8'h04;
      17'd9599: data = 8'h02;
      17'd9600: data = 8'h02;
      17'd9601: data = 8'h02;
      17'd9602: data = 8'h01;
      17'd9603: data = 8'h05;
      17'd9604: data = 8'h09;
      17'd9605: data = 8'h0a;
      17'd9606: data = 8'h05;
      17'd9607: data = 8'h05;
      17'd9608: data = 8'h05;
      17'd9609: data = 8'h06;
      17'd9610: data = 8'h0a;
      17'd9611: data = 8'h04;
      17'd9612: data = 8'h00;
      17'd9613: data = 8'h06;
      17'd9614: data = 8'h0e;
      17'd9615: data = 8'h0a;
      17'd9616: data = 8'h05;
      17'd9617: data = 8'h05;
      17'd9618: data = 8'h09;
      17'd9619: data = 8'h06;
      17'd9620: data = 8'h06;
      17'd9621: data = 8'h09;
      17'd9622: data = 8'h0d;
      17'd9623: data = 8'h11;
      17'd9624: data = 8'h0a;
      17'd9625: data = 8'hfe;
      17'd9626: data = 8'hf4;
      17'd9627: data = 8'hfe;
      17'd9628: data = 8'h05;
      17'd9629: data = 8'h06;
      17'd9630: data = 8'h0a;
      17'd9631: data = 8'h13;
      17'd9632: data = 8'h0e;
      17'd9633: data = 8'h00;
      17'd9634: data = 8'hfd;
      17'd9635: data = 8'hfd;
      17'd9636: data = 8'h00;
      17'd9637: data = 8'h05;
      17'd9638: data = 8'h0a;
      17'd9639: data = 8'h05;
      17'd9640: data = 8'hfe;
      17'd9641: data = 8'hf9;
      17'd9642: data = 8'hf4;
      17'd9643: data = 8'hf4;
      17'd9644: data = 8'h02;
      17'd9645: data = 8'h0a;
      17'd9646: data = 8'h01;
      17'd9647: data = 8'hf9;
      17'd9648: data = 8'hef;
      17'd9649: data = 8'hf1;
      17'd9650: data = 8'hf1;
      17'd9651: data = 8'hf4;
      17'd9652: data = 8'hf9;
      17'd9653: data = 8'hfe;
      17'd9654: data = 8'hfc;
      17'd9655: data = 8'he7;
      17'd9656: data = 8'he2;
      17'd9657: data = 8'hec;
      17'd9658: data = 8'hf1;
      17'd9659: data = 8'hec;
      17'd9660: data = 8'he7;
      17'd9661: data = 8'hed;
      17'd9662: data = 8'hf1;
      17'd9663: data = 8'he7;
      17'd9664: data = 8'he5;
      17'd9665: data = 8'he2;
      17'd9666: data = 8'he3;
      17'd9667: data = 8'hec;
      17'd9668: data = 8'heb;
      17'd9669: data = 8'heb;
      17'd9670: data = 8'he2;
      17'd9671: data = 8'hda;
      17'd9672: data = 8'he0;
      17'd9673: data = 8'hdb;
      17'd9674: data = 8'he4;
      17'd9675: data = 8'hed;
      17'd9676: data = 8'he9;
      17'd9677: data = 8'hda;
      17'd9678: data = 8'hde;
      17'd9679: data = 8'he7;
      17'd9680: data = 8'he0;
      17'd9681: data = 8'hde;
      17'd9682: data = 8'he5;
      17'd9683: data = 8'hf2;
      17'd9684: data = 8'hec;
      17'd9685: data = 8'hf1;
      17'd9686: data = 8'heb;
      17'd9687: data = 8'he4;
      17'd9688: data = 8'hf5;
      17'd9689: data = 8'hf4;
      17'd9690: data = 8'hf2;
      17'd9691: data = 8'hf2;
      17'd9692: data = 8'h01;
      17'd9693: data = 8'h01;
      17'd9694: data = 8'he5;
      17'd9695: data = 8'h01;
      17'd9696: data = 8'h19;
      17'd9697: data = 8'h19;
      17'd9698: data = 8'h05;
      17'd9699: data = 8'h04;
      17'd9700: data = 8'h15;
      17'd9701: data = 8'h06;
      17'd9702: data = 8'h0d;
      17'd9703: data = 8'h1e;
      17'd9704: data = 8'h22;
      17'd9705: data = 8'h12;
      17'd9706: data = 8'h12;
      17'd9707: data = 8'h13;
      17'd9708: data = 8'h11;
      17'd9709: data = 8'h1a;
      17'd9710: data = 8'h29;
      17'd9711: data = 8'h26;
      17'd9712: data = 8'h13;
      17'd9713: data = 8'h27;
      17'd9714: data = 8'h2c;
      17'd9715: data = 8'h1b;
      17'd9716: data = 8'h15;
      17'd9717: data = 8'h13;
      17'd9718: data = 8'h1c;
      17'd9719: data = 8'h1a;
      17'd9720: data = 8'h2b;
      17'd9721: data = 8'h33;
      17'd9722: data = 8'h16;
      17'd9723: data = 8'h05;
      17'd9724: data = 8'h0a;
      17'd9725: data = 8'h12;
      17'd9726: data = 8'h0e;
      17'd9727: data = 8'h26;
      17'd9728: data = 8'h2c;
      17'd9729: data = 8'h15;
      17'd9730: data = 8'h0d;
      17'd9731: data = 8'h04;
      17'd9732: data = 8'h00;
      17'd9733: data = 8'h05;
      17'd9734: data = 8'h12;
      17'd9735: data = 8'h16;
      17'd9736: data = 8'h09;
      17'd9737: data = 8'h02;
      17'd9738: data = 8'h00;
      17'd9739: data = 8'hfc;
      17'd9740: data = 8'hf9;
      17'd9741: data = 8'h01;
      17'd9742: data = 8'h0a;
      17'd9743: data = 8'hfc;
      17'd9744: data = 8'hed;
      17'd9745: data = 8'hfe;
      17'd9746: data = 8'h01;
      17'd9747: data = 8'hef;
      17'd9748: data = 8'hfc;
      17'd9749: data = 8'h01;
      17'd9750: data = 8'hf5;
      17'd9751: data = 8'hed;
      17'd9752: data = 8'hed;
      17'd9753: data = 8'hf2;
      17'd9754: data = 8'hf1;
      17'd9755: data = 8'h05;
      17'd9756: data = 8'h09;
      17'd9757: data = 8'hfc;
      17'd9758: data = 8'hf2;
      17'd9759: data = 8'heb;
      17'd9760: data = 8'heb;
      17'd9761: data = 8'heb;
      17'd9762: data = 8'h00;
      17'd9763: data = 8'h12;
      17'd9764: data = 8'h11;
      17'd9765: data = 8'hfc;
      17'd9766: data = 8'hef;
      17'd9767: data = 8'hef;
      17'd9768: data = 8'hf2;
      17'd9769: data = 8'h01;
      17'd9770: data = 8'h15;
      17'd9771: data = 8'h1c;
      17'd9772: data = 8'h04;
      17'd9773: data = 8'hf2;
      17'd9774: data = 8'hec;
      17'd9775: data = 8'hf2;
      17'd9776: data = 8'h05;
      17'd9777: data = 8'h19;
      17'd9778: data = 8'h23;
      17'd9779: data = 8'h15;
      17'd9780: data = 8'h04;
      17'd9781: data = 8'hfe;
      17'd9782: data = 8'hf6;
      17'd9783: data = 8'hfc;
      17'd9784: data = 8'h0e;
      17'd9785: data = 8'h1c;
      17'd9786: data = 8'h1b;
      17'd9787: data = 8'h11;
      17'd9788: data = 8'h05;
      17'd9789: data = 8'hfa;
      17'd9790: data = 8'hf6;
      17'd9791: data = 8'hfe;
      17'd9792: data = 8'h12;
      17'd9793: data = 8'h1c;
      17'd9794: data = 8'h13;
      17'd9795: data = 8'h01;
      17'd9796: data = 8'hf9;
      17'd9797: data = 8'hf5;
      17'd9798: data = 8'hf5;
      17'd9799: data = 8'h04;
      17'd9800: data = 8'h0e;
      17'd9801: data = 8'h0a;
      17'd9802: data = 8'h04;
      17'd9803: data = 8'hfc;
      17'd9804: data = 8'hef;
      17'd9805: data = 8'hed;
      17'd9806: data = 8'hf6;
      17'd9807: data = 8'h04;
      17'd9808: data = 8'h04;
      17'd9809: data = 8'hfd;
      17'd9810: data = 8'hf6;
      17'd9811: data = 8'hf4;
      17'd9812: data = 8'hf4;
      17'd9813: data = 8'hf2;
      17'd9814: data = 8'hf9;
      17'd9815: data = 8'hfe;
      17'd9816: data = 8'hf6;
      17'd9817: data = 8'hf5;
      17'd9818: data = 8'hf5;
      17'd9819: data = 8'hf1;
      17'd9820: data = 8'hef;
      17'd9821: data = 8'hf5;
      17'd9822: data = 8'hfe;
      17'd9823: data = 8'hfc;
      17'd9824: data = 8'hfd;
      17'd9825: data = 8'hfd;
      17'd9826: data = 8'hf9;
      17'd9827: data = 8'hf5;
      17'd9828: data = 8'hfa;
      17'd9829: data = 8'hfe;
      17'd9830: data = 8'hfa;
      17'd9831: data = 8'hfa;
      17'd9832: data = 8'hfd;
      17'd9833: data = 8'hfc;
      17'd9834: data = 8'hfc;
      17'd9835: data = 8'hfd;
      17'd9836: data = 8'h00;
      17'd9837: data = 8'h02;
      17'd9838: data = 8'h00;
      17'd9839: data = 8'hfe;
      17'd9840: data = 8'hfe;
      17'd9841: data = 8'hfd;
      17'd9842: data = 8'h01;
      17'd9843: data = 8'h05;
      17'd9844: data = 8'h02;
      17'd9845: data = 8'h01;
      17'd9846: data = 8'hfe;
      17'd9847: data = 8'hfe;
      17'd9848: data = 8'h01;
      17'd9849: data = 8'h02;
      17'd9850: data = 8'h05;
      17'd9851: data = 8'h04;
      17'd9852: data = 8'h01;
      17'd9853: data = 8'h02;
      17'd9854: data = 8'h04;
      17'd9855: data = 8'h04;
      17'd9856: data = 8'h04;
      17'd9857: data = 8'h06;
      17'd9858: data = 8'h0a;
      17'd9859: data = 8'h02;
      17'd9860: data = 8'hfa;
      17'd9861: data = 8'h00;
      17'd9862: data = 8'h02;
      17'd9863: data = 8'h02;
      17'd9864: data = 8'h05;
      17'd9865: data = 8'h0c;
      17'd9866: data = 8'h05;
      17'd9867: data = 8'hfd;
      17'd9868: data = 8'hfc;
      17'd9869: data = 8'hfc;
      17'd9870: data = 8'hfe;
      17'd9871: data = 8'h02;
      17'd9872: data = 8'h09;
      17'd9873: data = 8'h0a;
      17'd9874: data = 8'h04;
      17'd9875: data = 8'hfc;
      17'd9876: data = 8'hf5;
      17'd9877: data = 8'hef;
      17'd9878: data = 8'hf2;
      17'd9879: data = 8'h00;
      17'd9880: data = 8'h04;
      17'd9881: data = 8'hfd;
      17'd9882: data = 8'hfa;
      17'd9883: data = 8'hf4;
      17'd9884: data = 8'hef;
      17'd9885: data = 8'hed;
      17'd9886: data = 8'hf5;
      17'd9887: data = 8'hfd;
      17'd9888: data = 8'hfd;
      17'd9889: data = 8'hf5;
      17'd9890: data = 8'he9;
      17'd9891: data = 8'he5;
      17'd9892: data = 8'he7;
      17'd9893: data = 8'heb;
      17'd9894: data = 8'hf5;
      17'd9895: data = 8'hf5;
      17'd9896: data = 8'hf2;
      17'd9897: data = 8'hed;
      17'd9898: data = 8'he5;
      17'd9899: data = 8'he2;
      17'd9900: data = 8'he3;
      17'd9901: data = 8'he9;
      17'd9902: data = 8'hed;
      17'd9903: data = 8'hed;
      17'd9904: data = 8'he9;
      17'd9905: data = 8'he9;
      17'd9906: data = 8'he5;
      17'd9907: data = 8'hdc;
      17'd9908: data = 8'hde;
      17'd9909: data = 8'he4;
      17'd9910: data = 8'he9;
      17'd9911: data = 8'he4;
      17'd9912: data = 8'he5;
      17'd9913: data = 8'he5;
      17'd9914: data = 8'he2;
      17'd9915: data = 8'he3;
      17'd9916: data = 8'hdc;
      17'd9917: data = 8'he2;
      17'd9918: data = 8'he5;
      17'd9919: data = 8'he7;
      17'd9920: data = 8'he9;
      17'd9921: data = 8'he9;
      17'd9922: data = 8'hec;
      17'd9923: data = 8'he7;
      17'd9924: data = 8'he3;
      17'd9925: data = 8'he4;
      17'd9926: data = 8'hec;
      17'd9927: data = 8'hed;
      17'd9928: data = 8'hf4;
      17'd9929: data = 8'h00;
      17'd9930: data = 8'hfe;
      17'd9931: data = 8'h05;
      17'd9932: data = 8'hfa;
      17'd9933: data = 8'heb;
      17'd9934: data = 8'hef;
      17'd9935: data = 8'h05;
      17'd9936: data = 8'h13;
      17'd9937: data = 8'h05;
      17'd9938: data = 8'h05;
      17'd9939: data = 8'h12;
      17'd9940: data = 8'h06;
      17'd9941: data = 8'hfe;
      17'd9942: data = 8'h11;
      17'd9943: data = 8'h11;
      17'd9944: data = 8'h0d;
      17'd9945: data = 8'h0d;
      17'd9946: data = 8'h1a;
      17'd9947: data = 8'h27;
      17'd9948: data = 8'h1c;
      17'd9949: data = 8'h16;
      17'd9950: data = 8'h11;
      17'd9951: data = 8'h0c;
      17'd9952: data = 8'h1f;
      17'd9953: data = 8'h23;
      17'd9954: data = 8'h19;
      17'd9955: data = 8'h19;
      17'd9956: data = 8'h1f;
      17'd9957: data = 8'h1f;
      17'd9958: data = 8'h11;
      17'd9959: data = 8'h19;
      17'd9960: data = 8'h22;
      17'd9961: data = 8'h1f;
      17'd9962: data = 8'h15;
      17'd9963: data = 8'h19;
      17'd9964: data = 8'h1b;
      17'd9965: data = 8'h13;
      17'd9966: data = 8'h11;
      17'd9967: data = 8'h0d;
      17'd9968: data = 8'h0d;
      17'd9969: data = 8'h0d;
      17'd9970: data = 8'h0e;
      17'd9971: data = 8'h16;
      17'd9972: data = 8'h13;
      17'd9973: data = 8'h01;
      17'd9974: data = 8'h01;
      17'd9975: data = 8'hfd;
      17'd9976: data = 8'h00;
      17'd9977: data = 8'h09;
      17'd9978: data = 8'h09;
      17'd9979: data = 8'h0c;
      17'd9980: data = 8'h01;
      17'd9981: data = 8'hfa;
      17'd9982: data = 8'hfc;
      17'd9983: data = 8'hfe;
      17'd9984: data = 8'hf4;
      17'd9985: data = 8'hec;
      17'd9986: data = 8'hfc;
      17'd9987: data = 8'h01;
      17'd9988: data = 8'hfe;
      17'd9989: data = 8'h02;
      17'd9990: data = 8'hf6;
      17'd9991: data = 8'hed;
      17'd9992: data = 8'hef;
      17'd9993: data = 8'hef;
      17'd9994: data = 8'hf6;
      17'd9995: data = 8'hfe;
      17'd9996: data = 8'h06;
      17'd9997: data = 8'h0a;
      17'd9998: data = 8'hfa;
      17'd9999: data = 8'hed;
      17'd10000: data = 8'he9;
      17'd10001: data = 8'he7;
      17'd10002: data = 8'hf9;
      17'd10003: data = 8'h0d;
      17'd10004: data = 8'h11;
      17'd10005: data = 8'h04;
      17'd10006: data = 8'h00;
      17'd10007: data = 8'hf4;
      17'd10008: data = 8'hec;
      17'd10009: data = 8'hfe;
      17'd10010: data = 8'h0c;
      17'd10011: data = 8'h15;
      17'd10012: data = 8'h19;
      17'd10013: data = 8'h0c;
      17'd10014: data = 8'hfd;
      17'd10015: data = 8'hf4;
      17'd10016: data = 8'hf4;
      17'd10017: data = 8'h05;
      17'd10018: data = 8'h1b;
      17'd10019: data = 8'h23;
      17'd10020: data = 8'h22;
      17'd10021: data = 8'h11;
      17'd10022: data = 8'hfa;
      17'd10023: data = 8'hfa;
      17'd10024: data = 8'h05;
      17'd10025: data = 8'h0e;
      17'd10026: data = 8'h16;
      17'd10027: data = 8'h1e;
      17'd10028: data = 8'h1b;
      17'd10029: data = 8'h0a;
      17'd10030: data = 8'hfe;
      17'd10031: data = 8'hfe;
      17'd10032: data = 8'h09;
      17'd10033: data = 8'h15;
      17'd10034: data = 8'h1a;
      17'd10035: data = 8'h15;
      17'd10036: data = 8'h06;
      17'd10037: data = 8'hf9;
      17'd10038: data = 8'hfc;
      17'd10039: data = 8'h01;
      17'd10040: data = 8'h04;
      17'd10041: data = 8'h0a;
      17'd10042: data = 8'h09;
      17'd10043: data = 8'h01;
      17'd10044: data = 8'hfd;
      17'd10045: data = 8'hfa;
      17'd10046: data = 8'hfa;
      17'd10047: data = 8'hf6;
      17'd10048: data = 8'hfe;
      17'd10049: data = 8'h01;
      17'd10050: data = 8'hfe;
      17'd10051: data = 8'hfa;
      17'd10052: data = 8'hf4;
      17'd10053: data = 8'hf9;
      17'd10054: data = 8'hf9;
      17'd10055: data = 8'hf9;
      17'd10056: data = 8'hfa;
      17'd10057: data = 8'hf9;
      17'd10058: data = 8'hf6;
      17'd10059: data = 8'hf5;
      17'd10060: data = 8'hf6;
      17'd10061: data = 8'hf6;
      17'd10062: data = 8'hfc;
      17'd10063: data = 8'hfd;
      17'd10064: data = 8'hfd;
      17'd10065: data = 8'hfa;
      17'd10066: data = 8'hfc;
      17'd10067: data = 8'hfc;
      17'd10068: data = 8'hfa;
      17'd10069: data = 8'hfe;
      17'd10070: data = 8'hfc;
      17'd10071: data = 8'hfa;
      17'd10072: data = 8'hfc;
      17'd10073: data = 8'hf6;
      17'd10074: data = 8'hf9;
      17'd10075: data = 8'h01;
      17'd10076: data = 8'h02;
      17'd10077: data = 8'h02;
      17'd10078: data = 8'h00;
      17'd10079: data = 8'hfd;
      17'd10080: data = 8'hfd;
      17'd10081: data = 8'h00;
      17'd10082: data = 8'h01;
      17'd10083: data = 8'h00;
      17'd10084: data = 8'h02;
      17'd10085: data = 8'h00;
      17'd10086: data = 8'hfe;
      17'd10087: data = 8'h01;
      17'd10088: data = 8'hfe;
      17'd10089: data = 8'hfe;
      17'd10090: data = 8'h05;
      17'd10091: data = 8'h05;
      17'd10092: data = 8'h04;
      17'd10093: data = 8'h04;
      17'd10094: data = 8'hfe;
      17'd10095: data = 8'hfe;
      17'd10096: data = 8'h02;
      17'd10097: data = 8'h04;
      17'd10098: data = 8'h02;
      17'd10099: data = 8'h00;
      17'd10100: data = 8'h01;
      17'd10101: data = 8'h02;
      17'd10102: data = 8'h04;
      17'd10103: data = 8'h05;
      17'd10104: data = 8'h06;
      17'd10105: data = 8'h04;
      17'd10106: data = 8'hfd;
      17'd10107: data = 8'hfc;
      17'd10108: data = 8'hf6;
      17'd10109: data = 8'hf9;
      17'd10110: data = 8'h02;
      17'd10111: data = 8'h06;
      17'd10112: data = 8'h06;
      17'd10113: data = 8'h0d;
      17'd10114: data = 8'h05;
      17'd10115: data = 8'hf4;
      17'd10116: data = 8'hf1;
      17'd10117: data = 8'hec;
      17'd10118: data = 8'hf5;
      17'd10119: data = 8'h05;
      17'd10120: data = 8'h0d;
      17'd10121: data = 8'h02;
      17'd10122: data = 8'hfc;
      17'd10123: data = 8'hfd;
      17'd10124: data = 8'hf2;
      17'd10125: data = 8'hec;
      17'd10126: data = 8'hf9;
      17'd10127: data = 8'h00;
      17'd10128: data = 8'hfe;
      17'd10129: data = 8'hfc;
      17'd10130: data = 8'hf4;
      17'd10131: data = 8'hed;
      17'd10132: data = 8'hef;
      17'd10133: data = 8'hf5;
      17'd10134: data = 8'hfa;
      17'd10135: data = 8'hfa;
      17'd10136: data = 8'hf6;
      17'd10137: data = 8'hef;
      17'd10138: data = 8'he9;
      17'd10139: data = 8'he5;
      17'd10140: data = 8'he9;
      17'd10141: data = 8'heb;
      17'd10142: data = 8'hf1;
      17'd10143: data = 8'hf2;
      17'd10144: data = 8'hf6;
      17'd10145: data = 8'hf6;
      17'd10146: data = 8'hed;
      17'd10147: data = 8'he5;
      17'd10148: data = 8'he5;
      17'd10149: data = 8'he9;
      17'd10150: data = 8'heb;
      17'd10151: data = 8'he7;
      17'd10152: data = 8'he4;
      17'd10153: data = 8'he4;
      17'd10154: data = 8'he7;
      17'd10155: data = 8'heb;
      17'd10156: data = 8'hef;
      17'd10157: data = 8'hed;
      17'd10158: data = 8'he7;
      17'd10159: data = 8'he7;
      17'd10160: data = 8'he5;
      17'd10161: data = 8'he5;
      17'd10162: data = 8'heb;
      17'd10163: data = 8'hec;
      17'd10164: data = 8'hef;
      17'd10165: data = 8'heb;
      17'd10166: data = 8'he3;
      17'd10167: data = 8'he5;
      17'd10168: data = 8'heb;
      17'd10169: data = 8'hf5;
      17'd10170: data = 8'hf4;
      17'd10171: data = 8'hec;
      17'd10172: data = 8'hf2;
      17'd10173: data = 8'hf4;
      17'd10174: data = 8'hf1;
      17'd10175: data = 8'hf2;
      17'd10176: data = 8'h00;
      17'd10177: data = 8'hfd;
      17'd10178: data = 8'h02;
      17'd10179: data = 8'h04;
      17'd10180: data = 8'h01;
      17'd10181: data = 8'h00;
      17'd10182: data = 8'hf1;
      17'd10183: data = 8'hfe;
      17'd10184: data = 8'h01;
      17'd10185: data = 8'h06;
      17'd10186: data = 8'h1f;
      17'd10187: data = 8'h1b;
      17'd10188: data = 8'h09;
      17'd10189: data = 8'h09;
      17'd10190: data = 8'h0e;
      17'd10191: data = 8'h0c;
      17'd10192: data = 8'h11;
      17'd10193: data = 8'h1f;
      17'd10194: data = 8'h22;
      17'd10195: data = 8'h1a;
      17'd10196: data = 8'h13;
      17'd10197: data = 8'h09;
      17'd10198: data = 8'h0d;
      17'd10199: data = 8'h1e;
      17'd10200: data = 8'h22;
      17'd10201: data = 8'h15;
      17'd10202: data = 8'h15;
      17'd10203: data = 8'h2b;
      17'd10204: data = 8'h24;
      17'd10205: data = 8'h11;
      17'd10206: data = 8'h11;
      17'd10207: data = 8'h0e;
      17'd10208: data = 8'h0d;
      17'd10209: data = 8'h12;
      17'd10210: data = 8'h1f;
      17'd10211: data = 8'h1c;
      17'd10212: data = 8'h15;
      17'd10213: data = 8'h16;
      17'd10214: data = 8'h06;
      17'd10215: data = 8'h02;
      17'd10216: data = 8'h15;
      17'd10217: data = 8'h15;
      17'd10218: data = 8'h01;
      17'd10219: data = 8'h01;
      17'd10220: data = 8'h19;
      17'd10221: data = 8'h0d;
      17'd10222: data = 8'hfa;
      17'd10223: data = 8'h00;
      17'd10224: data = 8'h05;
      17'd10225: data = 8'h04;
      17'd10226: data = 8'h00;
      17'd10227: data = 8'hfd;
      17'd10228: data = 8'hf5;
      17'd10229: data = 8'hfc;
      17'd10230: data = 8'h04;
      17'd10231: data = 8'hfa;
      17'd10232: data = 8'hf5;
      17'd10233: data = 8'hfd;
      17'd10234: data = 8'hfc;
      17'd10235: data = 8'hef;
      17'd10236: data = 8'hf4;
      17'd10237: data = 8'hfd;
      17'd10238: data = 8'hfd;
      17'd10239: data = 8'h09;
      17'd10240: data = 8'h05;
      17'd10241: data = 8'hf4;
      17'd10242: data = 8'hed;
      17'd10243: data = 8'hed;
      17'd10244: data = 8'hed;
      17'd10245: data = 8'hfd;
      17'd10246: data = 8'h13;
      17'd10247: data = 8'h12;
      17'd10248: data = 8'h05;
      17'd10249: data = 8'hfc;
      17'd10250: data = 8'he7;
      17'd10251: data = 8'hed;
      17'd10252: data = 8'h09;
      17'd10253: data = 8'h09;
      17'd10254: data = 8'h0e;
      17'd10255: data = 8'h1a;
      17'd10256: data = 8'h0d;
      17'd10257: data = 8'hfa;
      17'd10258: data = 8'hf1;
      17'd10259: data = 8'h00;
      17'd10260: data = 8'h15;
      17'd10261: data = 8'h23;
      17'd10262: data = 8'h23;
      17'd10263: data = 8'h15;
      17'd10264: data = 8'h01;
      17'd10265: data = 8'hfa;
      17'd10266: data = 8'hfe;
      17'd10267: data = 8'h05;
      17'd10268: data = 8'h16;
      17'd10269: data = 8'h26;
      17'd10270: data = 8'h1f;
      17'd10271: data = 8'h0e;
      17'd10272: data = 8'h02;
      17'd10273: data = 8'hfe;
      17'd10274: data = 8'h04;
      17'd10275: data = 8'h0a;
      17'd10276: data = 8'h11;
      17'd10277: data = 8'h16;
      17'd10278: data = 8'h12;
      17'd10279: data = 8'hfe;
      17'd10280: data = 8'hf1;
      17'd10281: data = 8'hf6;
      17'd10282: data = 8'h04;
      17'd10283: data = 8'h0c;
      17'd10284: data = 8'h0c;
      17'd10285: data = 8'h04;
      17'd10286: data = 8'hfd;
      17'd10287: data = 8'hf5;
      17'd10288: data = 8'hf1;
      17'd10289: data = 8'hf1;
      17'd10290: data = 8'hf4;
      17'd10291: data = 8'h00;
      17'd10292: data = 8'h02;
      17'd10293: data = 8'hf9;
      17'd10294: data = 8'hf1;
      17'd10295: data = 8'hf4;
      17'd10296: data = 8'hf5;
      17'd10297: data = 8'hf1;
      17'd10298: data = 8'hf5;
      17'd10299: data = 8'hfc;
      17'd10300: data = 8'hf5;
      17'd10301: data = 8'hf2;
      17'd10302: data = 8'hf4;
      17'd10303: data = 8'hf2;
      17'd10304: data = 8'hf6;
      17'd10305: data = 8'hfa;
      17'd10306: data = 8'hfa;
      17'd10307: data = 8'hf5;
      17'd10308: data = 8'hf9;
      17'd10309: data = 8'hfc;
      17'd10310: data = 8'hf5;
      17'd10311: data = 8'hf6;
      17'd10312: data = 8'hf9;
      17'd10313: data = 8'hfc;
      17'd10314: data = 8'hfd;
      17'd10315: data = 8'hf9;
      17'd10316: data = 8'hf6;
      17'd10317: data = 8'hfe;
      17'd10318: data = 8'h01;
      17'd10319: data = 8'hfd;
      17'd10320: data = 8'hfd;
      17'd10321: data = 8'h00;
      17'd10322: data = 8'hfe;
      17'd10323: data = 8'hf9;
      17'd10324: data = 8'hfd;
      17'd10325: data = 8'hfe;
      17'd10326: data = 8'h01;
      17'd10327: data = 8'h02;
      17'd10328: data = 8'h04;
      17'd10329: data = 8'h02;
      17'd10330: data = 8'hfe;
      17'd10331: data = 8'h01;
      17'd10332: data = 8'h01;
      17'd10333: data = 8'hfe;
      17'd10334: data = 8'h00;
      17'd10335: data = 8'h05;
      17'd10336: data = 8'h05;
      17'd10337: data = 8'h00;
      17'd10338: data = 8'h01;
      17'd10339: data = 8'h04;
      17'd10340: data = 8'h06;
      17'd10341: data = 8'h0a;
      17'd10342: data = 8'h02;
      17'd10343: data = 8'h01;
      17'd10344: data = 8'h05;
      17'd10345: data = 8'h02;
      17'd10346: data = 8'h01;
      17'd10347: data = 8'h00;
      17'd10348: data = 8'h01;
      17'd10349: data = 8'h06;
      17'd10350: data = 8'h05;
      17'd10351: data = 8'h01;
      17'd10352: data = 8'h04;
      17'd10353: data = 8'h05;
      17'd10354: data = 8'h02;
      17'd10355: data = 8'h01;
      17'd10356: data = 8'h02;
      17'd10357: data = 8'h04;
      17'd10358: data = 8'h02;
      17'd10359: data = 8'hfe;
      17'd10360: data = 8'hf9;
      17'd10361: data = 8'hfc;
      17'd10362: data = 8'hfe;
      17'd10363: data = 8'hfc;
      17'd10364: data = 8'hf6;
      17'd10365: data = 8'hfe;
      17'd10366: data = 8'h05;
      17'd10367: data = 8'hfe;
      17'd10368: data = 8'hf4;
      17'd10369: data = 8'hf9;
      17'd10370: data = 8'hfa;
      17'd10371: data = 8'hfa;
      17'd10372: data = 8'hf6;
      17'd10373: data = 8'hf1;
      17'd10374: data = 8'hf1;
      17'd10375: data = 8'hf6;
      17'd10376: data = 8'hf9;
      17'd10377: data = 8'hf2;
      17'd10378: data = 8'hef;
      17'd10379: data = 8'hef;
      17'd10380: data = 8'hed;
      17'd10381: data = 8'heb;
      17'd10382: data = 8'hec;
      17'd10383: data = 8'hf4;
      17'd10384: data = 8'hf2;
      17'd10385: data = 8'hec;
      17'd10386: data = 8'hec;
      17'd10387: data = 8'hed;
      17'd10388: data = 8'hef;
      17'd10389: data = 8'he9;
      17'd10390: data = 8'he4;
      17'd10391: data = 8'he5;
      17'd10392: data = 8'he9;
      17'd10393: data = 8'heb;
      17'd10394: data = 8'he2;
      17'd10395: data = 8'he2;
      17'd10396: data = 8'he9;
      17'd10397: data = 8'he9;
      17'd10398: data = 8'he5;
      17'd10399: data = 8'he5;
      17'd10400: data = 8'he5;
      17'd10401: data = 8'he4;
      17'd10402: data = 8'hec;
      17'd10403: data = 8'he9;
      17'd10404: data = 8'he5;
      17'd10405: data = 8'he7;
      17'd10406: data = 8'hec;
      17'd10407: data = 8'hf1;
      17'd10408: data = 8'he4;
      17'd10409: data = 8'he5;
      17'd10410: data = 8'hec;
      17'd10411: data = 8'hec;
      17'd10412: data = 8'hed;
      17'd10413: data = 8'hf9;
      17'd10414: data = 8'hfc;
      17'd10415: data = 8'hf4;
      17'd10416: data = 8'hec;
      17'd10417: data = 8'hed;
      17'd10418: data = 8'hfa;
      17'd10419: data = 8'h00;
      17'd10420: data = 8'h04;
      17'd10421: data = 8'h00;
      17'd10422: data = 8'h01;
      17'd10423: data = 8'h04;
      17'd10424: data = 8'h05;
      17'd10425: data = 8'h09;
      17'd10426: data = 8'hfd;
      17'd10427: data = 8'h0a;
      17'd10428: data = 8'h19;
      17'd10429: data = 8'h13;
      17'd10430: data = 8'h0e;
      17'd10431: data = 8'h12;
      17'd10432: data = 8'h13;
      17'd10433: data = 8'h12;
      17'd10434: data = 8'h13;
      17'd10435: data = 8'h1e;
      17'd10436: data = 8'h24;
      17'd10437: data = 8'h22;
      17'd10438: data = 8'h16;
      17'd10439: data = 8'h0d;
      17'd10440: data = 8'h16;
      17'd10441: data = 8'h1c;
      17'd10442: data = 8'h1b;
      17'd10443: data = 8'h1f;
      17'd10444: data = 8'h2b;
      17'd10445: data = 8'h22;
      17'd10446: data = 8'h1b;
      17'd10447: data = 8'h15;
      17'd10448: data = 8'h13;
      17'd10449: data = 8'h1f;
      17'd10450: data = 8'h27;
      17'd10451: data = 8'h22;
      17'd10452: data = 8'h0d;
      17'd10453: data = 8'h0e;
      17'd10454: data = 8'h15;
      17'd10455: data = 8'h1a;
      17'd10456: data = 8'h1a;
      17'd10457: data = 8'h0d;
      17'd10458: data = 8'h04;
      17'd10459: data = 8'h0a;
      17'd10460: data = 8'h12;
      17'd10461: data = 8'h13;
      17'd10462: data = 8'h11;
      17'd10463: data = 8'h05;
      17'd10464: data = 8'h02;
      17'd10465: data = 8'h0c;
      17'd10466: data = 8'h11;
      17'd10467: data = 8'h02;
      17'd10468: data = 8'hf5;
      17'd10469: data = 8'hfd;
      17'd10470: data = 8'hf4;
      17'd10471: data = 8'hf6;
      17'd10472: data = 8'h09;
      17'd10473: data = 8'h06;
      17'd10474: data = 8'hf4;
      17'd10475: data = 8'he9;
      17'd10476: data = 8'hec;
      17'd10477: data = 8'hf9;
      17'd10478: data = 8'h02;
      17'd10479: data = 8'h05;
      17'd10480: data = 8'h01;
      17'd10481: data = 8'h01;
      17'd10482: data = 8'hfc;
      17'd10483: data = 8'he5;
      17'd10484: data = 8'he4;
      17'd10485: data = 8'hf2;
      17'd10486: data = 8'hfd;
      17'd10487: data = 8'h01;
      17'd10488: data = 8'h01;
      17'd10489: data = 8'h01;
      17'd10490: data = 8'hfd;
      17'd10491: data = 8'h01;
      17'd10492: data = 8'hfe;
      17'd10493: data = 8'hf1;
      17'd10494: data = 8'hfa;
      17'd10495: data = 8'h12;
      17'd10496: data = 8'h0d;
      17'd10497: data = 8'h0c;
      17'd10498: data = 8'h12;
      17'd10499: data = 8'h02;
      17'd10500: data = 8'hf4;
      17'd10501: data = 8'hfd;
      17'd10502: data = 8'h0e;
      17'd10503: data = 8'h19;
      17'd10504: data = 8'h1c;
      17'd10505: data = 8'h16;
      17'd10506: data = 8'h04;
      17'd10507: data = 8'h00;
      17'd10508: data = 8'h09;
      17'd10509: data = 8'h11;
      17'd10510: data = 8'h0e;
      17'd10511: data = 8'h12;
      17'd10512: data = 8'h1b;
      17'd10513: data = 8'h1a;
      17'd10514: data = 8'h09;
      17'd10515: data = 8'hfe;
      17'd10516: data = 8'h01;
      17'd10517: data = 8'h05;
      17'd10518: data = 8'h06;
      17'd10519: data = 8'h11;
      17'd10520: data = 8'h11;
      17'd10521: data = 8'h06;
      17'd10522: data = 8'h00;
      17'd10523: data = 8'h04;
      17'd10524: data = 8'h01;
      17'd10525: data = 8'hfe;
      17'd10526: data = 8'h0a;
      17'd10527: data = 8'h0a;
      17'd10528: data = 8'hfc;
      17'd10529: data = 8'hf2;
      17'd10530: data = 8'hf2;
      17'd10531: data = 8'hed;
      17'd10532: data = 8'hf1;
      17'd10533: data = 8'hfd;
      17'd10534: data = 8'h04;
      17'd10535: data = 8'hfd;
      17'd10536: data = 8'hf1;
      17'd10537: data = 8'hec;
      17'd10538: data = 8'hf4;
      17'd10539: data = 8'hfd;
      17'd10540: data = 8'hfc;
      17'd10541: data = 8'hf9;
      17'd10542: data = 8'hf2;
      17'd10543: data = 8'hf1;
      17'd10544: data = 8'hf2;
      17'd10545: data = 8'hf4;
      17'd10546: data = 8'hf2;
      17'd10547: data = 8'hf6;
      17'd10548: data = 8'h00;
      17'd10549: data = 8'h00;
      17'd10550: data = 8'hf9;
      17'd10551: data = 8'hf4;
      17'd10552: data = 8'hf6;
      17'd10553: data = 8'hf9;
      17'd10554: data = 8'hfc;
      17'd10555: data = 8'h00;
      17'd10556: data = 8'h02;
      17'd10557: data = 8'h02;
      17'd10558: data = 8'hfd;
      17'd10559: data = 8'hf9;
      17'd10560: data = 8'hfd;
      17'd10561: data = 8'h04;
      17'd10562: data = 8'h02;
      17'd10563: data = 8'hfe;
      17'd10564: data = 8'h00;
      17'd10565: data = 8'h01;
      17'd10566: data = 8'h00;
      17'd10567: data = 8'hfd;
      17'd10568: data = 8'hfe;
      17'd10569: data = 8'h05;
      17'd10570: data = 8'h0d;
      17'd10571: data = 8'h0a;
      17'd10572: data = 8'h02;
      17'd10573: data = 8'h00;
      17'd10574: data = 8'h00;
      17'd10575: data = 8'h01;
      17'd10576: data = 8'h01;
      17'd10577: data = 8'h01;
      17'd10578: data = 8'h02;
      17'd10579: data = 8'h02;
      17'd10580: data = 8'h02;
      17'd10581: data = 8'h01;
      17'd10582: data = 8'h04;
      17'd10583: data = 8'h06;
      17'd10584: data = 8'h04;
      17'd10585: data = 8'h05;
      17'd10586: data = 8'h04;
      17'd10587: data = 8'h01;
      17'd10588: data = 8'hfe;
      17'd10589: data = 8'hfe;
      17'd10590: data = 8'h00;
      17'd10591: data = 8'h00;
      17'd10592: data = 8'h04;
      17'd10593: data = 8'h05;
      17'd10594: data = 8'hfd;
      17'd10595: data = 8'hfd;
      17'd10596: data = 8'h01;
      17'd10597: data = 8'h02;
      17'd10598: data = 8'hfd;
      17'd10599: data = 8'hfc;
      17'd10600: data = 8'h02;
      17'd10601: data = 8'h00;
      17'd10602: data = 8'hfd;
      17'd10603: data = 8'h02;
      17'd10604: data = 8'hfd;
      17'd10605: data = 8'hf5;
      17'd10606: data = 8'hf4;
      17'd10607: data = 8'hf1;
      17'd10608: data = 8'hf4;
      17'd10609: data = 8'hf5;
      17'd10610: data = 8'hf9;
      17'd10611: data = 8'hfc;
      17'd10612: data = 8'hfa;
      17'd10613: data = 8'hf9;
      17'd10614: data = 8'hf5;
      17'd10615: data = 8'hf2;
      17'd10616: data = 8'hed;
      17'd10617: data = 8'hed;
      17'd10618: data = 8'hf4;
      17'd10619: data = 8'hf2;
      17'd10620: data = 8'heb;
      17'd10621: data = 8'heb;
      17'd10622: data = 8'hed;
      17'd10623: data = 8'hed;
      17'd10624: data = 8'heb;
      17'd10625: data = 8'heb;
      17'd10626: data = 8'hec;
      17'd10627: data = 8'heb;
      17'd10628: data = 8'heb;
      17'd10629: data = 8'he9;
      17'd10630: data = 8'he7;
      17'd10631: data = 8'he5;
      17'd10632: data = 8'he5;
      17'd10633: data = 8'hed;
      17'd10634: data = 8'hed;
      17'd10635: data = 8'he7;
      17'd10636: data = 8'he7;
      17'd10637: data = 8'he5;
      17'd10638: data = 8'he4;
      17'd10639: data = 8'he5;
      17'd10640: data = 8'heb;
      17'd10641: data = 8'he9;
      17'd10642: data = 8'he3;
      17'd10643: data = 8'he3;
      17'd10644: data = 8'he9;
      17'd10645: data = 8'heb;
      17'd10646: data = 8'heb;
      17'd10647: data = 8'hf1;
      17'd10648: data = 8'hf6;
      17'd10649: data = 8'hec;
      17'd10650: data = 8'he9;
      17'd10651: data = 8'hef;
      17'd10652: data = 8'hed;
      17'd10653: data = 8'hf5;
      17'd10654: data = 8'hf6;
      17'd10655: data = 8'hf5;
      17'd10656: data = 8'hf4;
      17'd10657: data = 8'hef;
      17'd10658: data = 8'hfc;
      17'd10659: data = 8'hfe;
      17'd10660: data = 8'hfc;
      17'd10661: data = 8'hfc;
      17'd10662: data = 8'h04;
      17'd10663: data = 8'h05;
      17'd10664: data = 8'h01;
      17'd10665: data = 8'h09;
      17'd10666: data = 8'h04;
      17'd10667: data = 8'h04;
      17'd10668: data = 8'h0e;
      17'd10669: data = 8'h0e;
      17'd10670: data = 8'h12;
      17'd10671: data = 8'h15;
      17'd10672: data = 8'h0e;
      17'd10673: data = 8'h0e;
      17'd10674: data = 8'h0a;
      17'd10675: data = 8'h13;
      17'd10676: data = 8'h16;
      17'd10677: data = 8'h0e;
      17'd10678: data = 8'h1b;
      17'd10679: data = 8'h1c;
      17'd10680: data = 8'h23;
      17'd10681: data = 8'h1e;
      17'd10682: data = 8'h12;
      17'd10683: data = 8'h1c;
      17'd10684: data = 8'h13;
      17'd10685: data = 8'h12;
      17'd10686: data = 8'h12;
      17'd10687: data = 8'h1f;
      17'd10688: data = 8'h2c;
      17'd10689: data = 8'h16;
      17'd10690: data = 8'h1b;
      17'd10691: data = 8'h1b;
      17'd10692: data = 8'h0d;
      17'd10693: data = 8'h15;
      17'd10694: data = 8'h0e;
      17'd10695: data = 8'h11;
      17'd10696: data = 8'h1f;
      17'd10697: data = 8'h1b;
      17'd10698: data = 8'h16;
      17'd10699: data = 8'h11;
      17'd10700: data = 8'h09;
      17'd10701: data = 8'h00;
      17'd10702: data = 8'h01;
      17'd10703: data = 8'h0d;
      17'd10704: data = 8'h0a;
      17'd10705: data = 8'h12;
      17'd10706: data = 8'h1e;
      17'd10707: data = 8'h0a;
      17'd10708: data = 8'hfc;
      17'd10709: data = 8'h01;
      17'd10710: data = 8'hfa;
      17'd10711: data = 8'hef;
      17'd10712: data = 8'hef;
      17'd10713: data = 8'h00;
      17'd10714: data = 8'h05;
      17'd10715: data = 8'hfe;
      17'd10716: data = 8'h04;
      17'd10717: data = 8'h06;
      17'd10718: data = 8'hfc;
      17'd10719: data = 8'heb;
      17'd10720: data = 8'hed;
      17'd10721: data = 8'hef;
      17'd10722: data = 8'hf9;
      17'd10723: data = 8'h0a;
      17'd10724: data = 8'h05;
      17'd10725: data = 8'hfc;
      17'd10726: data = 8'hf5;
      17'd10727: data = 8'hf1;
      17'd10728: data = 8'hef;
      17'd10729: data = 8'hfc;
      17'd10730: data = 8'h0d;
      17'd10731: data = 8'h0e;
      17'd10732: data = 8'h09;
      17'd10733: data = 8'hfe;
      17'd10734: data = 8'hf9;
      17'd10735: data = 8'hf6;
      17'd10736: data = 8'hf9;
      17'd10737: data = 8'h01;
      17'd10738: data = 8'h0d;
      17'd10739: data = 8'h15;
      17'd10740: data = 8'h13;
      17'd10741: data = 8'h0c;
      17'd10742: data = 8'h01;
      17'd10743: data = 8'h02;
      17'd10744: data = 8'h0c;
      17'd10745: data = 8'h0e;
      17'd10746: data = 8'h12;
      17'd10747: data = 8'h13;
      17'd10748: data = 8'h11;
      17'd10749: data = 8'h06;
      17'd10750: data = 8'h0c;
      17'd10751: data = 8'h11;
      17'd10752: data = 8'h12;
      17'd10753: data = 8'h1a;
      17'd10754: data = 8'h1a;
      17'd10755: data = 8'h0d;
      17'd10756: data = 8'h04;
      17'd10757: data = 8'h01;
      17'd10758: data = 8'h02;
      17'd10759: data = 8'h0e;
      17'd10760: data = 8'h13;
      17'd10761: data = 8'h11;
      17'd10762: data = 8'h0c;
      17'd10763: data = 8'h04;
      17'd10764: data = 8'hfe;
      17'd10765: data = 8'h04;
      17'd10766: data = 8'h09;
      17'd10767: data = 8'h06;
      17'd10768: data = 8'h02;
      17'd10769: data = 8'hfc;
      17'd10770: data = 8'hf4;
      17'd10771: data = 8'hf1;
      17'd10772: data = 8'hf4;
      17'd10773: data = 8'hf5;
      17'd10774: data = 8'hfc;
      17'd10775: data = 8'h01;
      17'd10776: data = 8'h01;
      17'd10777: data = 8'hfa;
      17'd10778: data = 8'hf2;
      17'd10779: data = 8'hf2;
      17'd10780: data = 8'hf1;
      17'd10781: data = 8'hf1;
      17'd10782: data = 8'hf4;
      17'd10783: data = 8'hf9;
      17'd10784: data = 8'hf6;
      17'd10785: data = 8'hf4;
      17'd10786: data = 8'hf4;
      17'd10787: data = 8'hf6;
      17'd10788: data = 8'hfa;
      17'd10789: data = 8'hfc;
      17'd10790: data = 8'hf9;
      17'd10791: data = 8'hf9;
      17'd10792: data = 8'hfa;
      17'd10793: data = 8'hf6;
      17'd10794: data = 8'hf6;
      17'd10795: data = 8'hfd;
      17'd10796: data = 8'hfe;
      17'd10797: data = 8'h00;
      17'd10798: data = 8'h01;
      17'd10799: data = 8'hfd;
      17'd10800: data = 8'hfc;
      17'd10801: data = 8'h02;
      17'd10802: data = 8'h06;
      17'd10803: data = 8'h02;
      17'd10804: data = 8'h01;
      17'd10805: data = 8'h00;
      17'd10806: data = 8'hfd;
      17'd10807: data = 8'h00;
      17'd10808: data = 8'h04;
      17'd10809: data = 8'h06;
      17'd10810: data = 8'h0a;
      17'd10811: data = 8'h0d;
      17'd10812: data = 8'h0c;
      17'd10813: data = 8'h0a;
      17'd10814: data = 8'h05;
      17'd10815: data = 8'hfe;
      17'd10816: data = 8'hfe;
      17'd10817: data = 8'h04;
      17'd10818: data = 8'h05;
      17'd10819: data = 8'h06;
      17'd10820: data = 8'h0a;
      17'd10821: data = 8'h05;
      17'd10822: data = 8'h06;
      17'd10823: data = 8'h0a;
      17'd10824: data = 8'h06;
      17'd10825: data = 8'h09;
      17'd10826: data = 8'h09;
      17'd10827: data = 8'h09;
      17'd10828: data = 8'h04;
      17'd10829: data = 8'hfa;
      17'd10830: data = 8'hf9;
      17'd10831: data = 8'h00;
      17'd10832: data = 8'h01;
      17'd10833: data = 8'h0a;
      17'd10834: data = 8'h0e;
      17'd10835: data = 8'h0c;
      17'd10836: data = 8'h01;
      17'd10837: data = 8'hfa;
      17'd10838: data = 8'hf5;
      17'd10839: data = 8'hf5;
      17'd10840: data = 8'hfd;
      17'd10841: data = 8'h01;
      17'd10842: data = 8'h02;
      17'd10843: data = 8'h05;
      17'd10844: data = 8'h01;
      17'd10845: data = 8'hf2;
      17'd10846: data = 8'heb;
      17'd10847: data = 8'heb;
      17'd10848: data = 8'hed;
      17'd10849: data = 8'hf1;
      17'd10850: data = 8'hf5;
      17'd10851: data = 8'hf6;
      17'd10852: data = 8'hf4;
      17'd10853: data = 8'hf4;
      17'd10854: data = 8'hf2;
      17'd10855: data = 8'heb;
      17'd10856: data = 8'heb;
      17'd10857: data = 8'hec;
      17'd10858: data = 8'he9;
      17'd10859: data = 8'he5;
      17'd10860: data = 8'he7;
      17'd10861: data = 8'he9;
      17'd10862: data = 8'he9;
      17'd10863: data = 8'heb;
      17'd10864: data = 8'heb;
      17'd10865: data = 8'he5;
      17'd10866: data = 8'he4;
      17'd10867: data = 8'he4;
      17'd10868: data = 8'he3;
      17'd10869: data = 8'he5;
      17'd10870: data = 8'he7;
      17'd10871: data = 8'he4;
      17'd10872: data = 8'he2;
      17'd10873: data = 8'he7;
      17'd10874: data = 8'he5;
      17'd10875: data = 8'he3;
      17'd10876: data = 8'he5;
      17'd10877: data = 8'he5;
      17'd10878: data = 8'he7;
      17'd10879: data = 8'he5;
      17'd10880: data = 8'he5;
      17'd10881: data = 8'he4;
      17'd10882: data = 8'he4;
      17'd10883: data = 8'he5;
      17'd10884: data = 8'he7;
      17'd10885: data = 8'he4;
      17'd10886: data = 8'he4;
      17'd10887: data = 8'hec;
      17'd10888: data = 8'hef;
      17'd10889: data = 8'hf4;
      17'd10890: data = 8'hf5;
      17'd10891: data = 8'hf2;
      17'd10892: data = 8'hed;
      17'd10893: data = 8'heb;
      17'd10894: data = 8'hed;
      17'd10895: data = 8'hf4;
      17'd10896: data = 8'hf9;
      17'd10897: data = 8'hfa;
      17'd10898: data = 8'hfd;
      17'd10899: data = 8'h04;
      17'd10900: data = 8'h01;
      17'd10901: data = 8'hfe;
      17'd10902: data = 8'hfd;
      17'd10903: data = 8'hfd;
      17'd10904: data = 8'h01;
      17'd10905: data = 8'h0a;
      17'd10906: data = 8'h12;
      17'd10907: data = 8'h11;
      17'd10908: data = 8'h0c;
      17'd10909: data = 8'h09;
      17'd10910: data = 8'h09;
      17'd10911: data = 8'h0c;
      17'd10912: data = 8'h13;
      17'd10913: data = 8'h1a;
      17'd10914: data = 8'h1a;
      17'd10915: data = 8'h19;
      17'd10916: data = 8'h16;
      17'd10917: data = 8'h15;
      17'd10918: data = 8'h11;
      17'd10919: data = 8'h13;
      17'd10920: data = 8'h1a;
      17'd10921: data = 8'h1b;
      17'd10922: data = 8'h1f;
      17'd10923: data = 8'h1a;
      17'd10924: data = 8'h19;
      17'd10925: data = 8'h1c;
      17'd10926: data = 8'h19;
      17'd10927: data = 8'h15;
      17'd10928: data = 8'h06;
      17'd10929: data = 8'h19;
      17'd10930: data = 8'h22;
      17'd10931: data = 8'h16;
      17'd10932: data = 8'h23;
      17'd10933: data = 8'h15;
      17'd10934: data = 8'h09;
      17'd10935: data = 8'h09;
      17'd10936: data = 8'h0e;
      17'd10937: data = 8'h15;
      17'd10938: data = 8'h0a;
      17'd10939: data = 8'h0a;
      17'd10940: data = 8'h13;
      17'd10941: data = 8'h04;
      17'd10942: data = 8'h09;
      17'd10943: data = 8'h15;
      17'd10944: data = 8'h00;
      17'd10945: data = 8'h00;
      17'd10946: data = 8'h01;
      17'd10947: data = 8'h05;
      17'd10948: data = 8'h05;
      17'd10949: data = 8'h09;
      17'd10950: data = 8'h0a;
      17'd10951: data = 8'hf2;
      17'd10952: data = 8'he4;
      17'd10953: data = 8'he9;
      17'd10954: data = 8'he7;
      17'd10955: data = 8'hec;
      17'd10956: data = 8'hfc;
      17'd10957: data = 8'h09;
      17'd10958: data = 8'h15;
      17'd10959: data = 8'h04;
      17'd10960: data = 8'hf4;
      17'd10961: data = 8'hf2;
      17'd10962: data = 8'hec;
      17'd10963: data = 8'hec;
      17'd10964: data = 8'hec;
      17'd10965: data = 8'hed;
      17'd10966: data = 8'hfd;
      17'd10967: data = 8'h05;
      17'd10968: data = 8'h02;
      17'd10969: data = 8'h09;
      17'd10970: data = 8'h0c;
      17'd10971: data = 8'h04;
      17'd10972: data = 8'h04;
      17'd10973: data = 8'h04;
      17'd10974: data = 8'hfc;
      17'd10975: data = 8'hf6;
      17'd10976: data = 8'hfc;
      17'd10977: data = 8'h02;
      17'd10978: data = 8'h11;
      17'd10979: data = 8'h24;
      17'd10980: data = 8'h1f;
      17'd10981: data = 8'h0a;
      17'd10982: data = 8'h09;
      17'd10983: data = 8'h06;
      17'd10984: data = 8'h0e;
      17'd10985: data = 8'h16;
      17'd10986: data = 8'h0e;
      17'd10987: data = 8'h1a;
      17'd10988: data = 8'h11;
      17'd10989: data = 8'h05;
      17'd10990: data = 8'h0a;
      17'd10991: data = 8'h0e;
      17'd10992: data = 8'h1b;
      17'd10993: data = 8'h22;
      17'd10994: data = 8'h24;
      17'd10995: data = 8'h16;
      17'd10996: data = 8'h05;
      17'd10997: data = 8'h04;
      17'd10998: data = 8'h01;
      17'd10999: data = 8'h02;
      17'd11000: data = 8'h06;
      17'd11001: data = 8'h06;
      17'd11002: data = 8'h0c;
      17'd11003: data = 8'h01;
      17'd11004: data = 8'h01;
      17'd11005: data = 8'h0a;
      17'd11006: data = 8'h04;
      17'd11007: data = 8'hfe;
      17'd11008: data = 8'hf9;
      17'd11009: data = 8'hf9;
      17'd11010: data = 8'hed;
      17'd11011: data = 8'he5;
      17'd11012: data = 8'he9;
      17'd11013: data = 8'hed;
      17'd11014: data = 8'hfe;
      17'd11015: data = 8'h05;
      17'd11016: data = 8'h00;
      17'd11017: data = 8'hf6;
      17'd11018: data = 8'hed;
      17'd11019: data = 8'heb;
      17'd11020: data = 8'heb;
      17'd11021: data = 8'he9;
      17'd11022: data = 8'hed;
      17'd11023: data = 8'hf4;
      17'd11024: data = 8'hf2;
      17'd11025: data = 8'hec;
      17'd11026: data = 8'hf1;
      17'd11027: data = 8'hfd;
      17'd11028: data = 8'hfe;
      17'd11029: data = 8'h00;
      17'd11030: data = 8'hfe;
      17'd11031: data = 8'hfd;
      17'd11032: data = 8'hf5;
      17'd11033: data = 8'hed;
      17'd11034: data = 8'hf4;
      17'd11035: data = 8'hf9;
      17'd11036: data = 8'h00;
      17'd11037: data = 8'h05;
      17'd11038: data = 8'h06;
      17'd11039: data = 8'h0a;
      17'd11040: data = 8'h09;
      17'd11041: data = 8'h0c;
      17'd11042: data = 8'h0c;
      17'd11043: data = 8'h05;
      17'd11044: data = 8'h09;
      17'd11045: data = 8'h04;
      17'd11046: data = 8'h02;
      17'd11047: data = 8'h06;
      17'd11048: data = 8'h09;
      17'd11049: data = 8'h11;
      17'd11050: data = 8'h16;
      17'd11051: data = 8'h16;
      17'd11052: data = 8'h16;
      17'd11053: data = 8'h11;
      17'd11054: data = 8'h0c;
      17'd11055: data = 8'h05;
      17'd11056: data = 8'h04;
      17'd11057: data = 8'h09;
      17'd11058: data = 8'h06;
      17'd11059: data = 8'h0a;
      17'd11060: data = 8'h09;
      17'd11061: data = 8'h0c;
      17'd11062: data = 8'h0e;
      17'd11063: data = 8'h11;
      17'd11064: data = 8'h15;
      17'd11065: data = 8'h0d;
      17'd11066: data = 8'h01;
      17'd11067: data = 8'hf6;
      17'd11068: data = 8'hf9;
      17'd11069: data = 8'hf9;
      17'd11070: data = 8'hf4;
      17'd11071: data = 8'h00;
      17'd11072: data = 8'h15;
      17'd11073: data = 8'h16;
      17'd11074: data = 8'h0c;
      17'd11075: data = 8'h01;
      17'd11076: data = 8'hf9;
      17'd11077: data = 8'hed;
      17'd11078: data = 8'heb;
      17'd11079: data = 8'hf2;
      17'd11080: data = 8'hf4;
      17'd11081: data = 8'hfa;
      17'd11082: data = 8'hf9;
      17'd11083: data = 8'hf1;
      17'd11084: data = 8'hf4;
      17'd11085: data = 8'hf5;
      17'd11086: data = 8'hf5;
      17'd11087: data = 8'hed;
      17'd11088: data = 8'hec;
      17'd11089: data = 8'hed;
      17'd11090: data = 8'he5;
      17'd11091: data = 8'he4;
      17'd11092: data = 8'hde;
      17'd11093: data = 8'hdc;
      17'd11094: data = 8'hec;
      17'd11095: data = 8'hed;
      17'd11096: data = 8'he3;
      17'd11097: data = 8'he3;
      17'd11098: data = 8'he5;
      17'd11099: data = 8'he7;
      17'd11100: data = 8'hdc;
      17'd11101: data = 8'hdc;
      17'd11102: data = 8'he3;
      17'd11103: data = 8'hdb;
      17'd11104: data = 8'hda;
      17'd11105: data = 8'hd8;
      17'd11106: data = 8'hda;
      17'd11107: data = 8'he0;
      17'd11108: data = 8'he7;
      17'd11109: data = 8'heb;
      17'd11110: data = 8'he4;
      17'd11111: data = 8'he5;
      17'd11112: data = 8'hde;
      17'd11113: data = 8'hd5;
      17'd11114: data = 8'hd5;
      17'd11115: data = 8'hdb;
      17'd11116: data = 8'he5;
      17'd11117: data = 8'he9;
      17'd11118: data = 8'he7;
      17'd11119: data = 8'he9;
      17'd11120: data = 8'hed;
      17'd11121: data = 8'hef;
      17'd11122: data = 8'hed;
      17'd11123: data = 8'hef;
      17'd11124: data = 8'hef;
      17'd11125: data = 8'hec;
      17'd11126: data = 8'hec;
      17'd11127: data = 8'hec;
      17'd11128: data = 8'hef;
      17'd11129: data = 8'hfa;
      17'd11130: data = 8'h00;
      17'd11131: data = 8'h01;
      17'd11132: data = 8'h02;
      17'd11133: data = 8'h01;
      17'd11134: data = 8'h02;
      17'd11135: data = 8'hfd;
      17'd11136: data = 8'hfd;
      17'd11137: data = 8'h02;
      17'd11138: data = 8'h09;
      17'd11139: data = 8'h0d;
      17'd11140: data = 8'h0a;
      17'd11141: data = 8'h0e;
      17'd11142: data = 8'h12;
      17'd11143: data = 8'h16;
      17'd11144: data = 8'h1a;
      17'd11145: data = 8'h11;
      17'd11146: data = 8'h13;
      17'd11147: data = 8'h15;
      17'd11148: data = 8'h0e;
      17'd11149: data = 8'h0e;
      17'd11150: data = 8'h11;
      17'd11151: data = 8'h1f;
      17'd11152: data = 8'h22;
      17'd11153: data = 8'h22;
      17'd11154: data = 8'h1e;
      17'd11155: data = 8'h0e;
      17'd11156: data = 8'h1a;
      17'd11157: data = 8'h1c;
      17'd11158: data = 8'h0d;
      17'd11159: data = 8'h11;
      17'd11160: data = 8'h13;
      17'd11161: data = 8'h1b;
      17'd11162: data = 8'h16;
      17'd11163: data = 8'h0c;
      17'd11164: data = 8'h1b;
      17'd11165: data = 8'h19;
      17'd11166: data = 8'h0d;
      17'd11167: data = 8'h13;
      17'd11168: data = 8'h11;
      17'd11169: data = 8'h11;
      17'd11170: data = 8'h04;
      17'd11171: data = 8'h01;
      17'd11172: data = 8'h0c;
      17'd11173: data = 8'h06;
      17'd11174: data = 8'h0c;
      17'd11175: data = 8'h04;
      17'd11176: data = 8'hf1;
      17'd11177: data = 8'h02;
      17'd11178: data = 8'h0c;
      17'd11179: data = 8'h01;
      17'd11180: data = 8'h09;
      17'd11181: data = 8'h0d;
      17'd11182: data = 8'h11;
      17'd11183: data = 8'h05;
      17'd11184: data = 8'hf5;
      17'd11185: data = 8'heb;
      17'd11186: data = 8'hd6;
      17'd11187: data = 8'he4;
      17'd11188: data = 8'hf2;
      17'd11189: data = 8'he4;
      17'd11190: data = 8'hef;
      17'd11191: data = 8'h05;
      17'd11192: data = 8'h11;
      17'd11193: data = 8'h12;
      17'd11194: data = 8'h0c;
      17'd11195: data = 8'h06;
      17'd11196: data = 8'hf4;
      17'd11197: data = 8'he4;
      17'd11198: data = 8'he4;
      17'd11199: data = 8'hdb;
      17'd11200: data = 8'heb;
      17'd11201: data = 8'h06;
      17'd11202: data = 8'h04;
      17'd11203: data = 8'h15;
      17'd11204: data = 8'h26;
      17'd11205: data = 8'h16;
      17'd11206: data = 8'h06;
      17'd11207: data = 8'hfe;
      17'd11208: data = 8'hf9;
      17'd11209: data = 8'hf6;
      17'd11210: data = 8'hf6;
      17'd11211: data = 8'h00;
      17'd11212: data = 8'h02;
      17'd11213: data = 8'h15;
      17'd11214: data = 8'h29;
      17'd11215: data = 8'h1f;
      17'd11216: data = 8'h1b;
      17'd11217: data = 8'h1e;
      17'd11218: data = 8'h1c;
      17'd11219: data = 8'h0e;
      17'd11220: data = 8'h01;
      17'd11221: data = 8'h04;
      17'd11222: data = 8'h0a;
      17'd11223: data = 8'h0d;
      17'd11224: data = 8'h19;
      17'd11225: data = 8'h1a;
      17'd11226: data = 8'h22;
      17'd11227: data = 8'h23;
      17'd11228: data = 8'h15;
      17'd11229: data = 8'h12;
      17'd11230: data = 8'h13;
      17'd11231: data = 8'h11;
      17'd11232: data = 8'h0a;
      17'd11233: data = 8'h05;
      17'd11234: data = 8'hfe;
      17'd11235: data = 8'hfc;
      17'd11236: data = 8'h01;
      17'd11237: data = 8'hfd;
      17'd11238: data = 8'hfa;
      17'd11239: data = 8'h09;
      17'd11240: data = 8'h13;
      17'd11241: data = 8'h09;
      17'd11242: data = 8'hfc;
      17'd11243: data = 8'hf4;
      17'd11244: data = 8'hed;
      17'd11245: data = 8'he5;
      17'd11246: data = 8'he3;
      17'd11247: data = 8'he5;
      17'd11248: data = 8'he9;
      17'd11249: data = 8'hec;
      17'd11250: data = 8'hf2;
      17'd11251: data = 8'hf5;
      17'd11252: data = 8'hf5;
      17'd11253: data = 8'hf9;
      17'd11254: data = 8'hf4;
      17'd11255: data = 8'hec;
      17'd11256: data = 8'he5;
      17'd11257: data = 8'he4;
      17'd11258: data = 8'he2;
      17'd11259: data = 8'he2;
      17'd11260: data = 8'he9;
      17'd11261: data = 8'hf9;
      17'd11262: data = 8'h05;
      17'd11263: data = 8'h09;
      17'd11264: data = 8'h01;
      17'd11265: data = 8'h02;
      17'd11266: data = 8'h04;
      17'd11267: data = 8'hfc;
      17'd11268: data = 8'hf5;
      17'd11269: data = 8'hf5;
      17'd11270: data = 8'hf5;
      17'd11271: data = 8'hfd;
      17'd11272: data = 8'h02;
      17'd11273: data = 8'h09;
      17'd11274: data = 8'h12;
      17'd11275: data = 8'h19;
      17'd11276: data = 8'h1c;
      17'd11277: data = 8'h15;
      17'd11278: data = 8'h15;
      17'd11279: data = 8'h11;
      17'd11280: data = 8'h09;
      17'd11281: data = 8'h09;
      17'd11282: data = 8'h09;
      17'd11283: data = 8'h0e;
      17'd11284: data = 8'h15;
      17'd11285: data = 8'h1b;
      17'd11286: data = 8'h19;
      17'd11287: data = 8'h1b;
      17'd11288: data = 8'h1f;
      17'd11289: data = 8'h1f;
      17'd11290: data = 8'h1a;
      17'd11291: data = 8'h12;
      17'd11292: data = 8'h12;
      17'd11293: data = 8'h0d;
      17'd11294: data = 8'h09;
      17'd11295: data = 8'h0d;
      17'd11296: data = 8'h0c;
      17'd11297: data = 8'h11;
      17'd11298: data = 8'h11;
      17'd11299: data = 8'h0d;
      17'd11300: data = 8'h12;
      17'd11301: data = 8'h06;
      17'd11302: data = 8'h00;
      17'd11303: data = 8'h06;
      17'd11304: data = 8'h0a;
      17'd11305: data = 8'h04;
      17'd11306: data = 8'hfe;
      17'd11307: data = 8'h00;
      17'd11308: data = 8'hfa;
      17'd11309: data = 8'hf4;
      17'd11310: data = 8'hf4;
      17'd11311: data = 8'hf2;
      17'd11312: data = 8'hf4;
      17'd11313: data = 8'hf6;
      17'd11314: data = 8'hf2;
      17'd11315: data = 8'hed;
      17'd11316: data = 8'he9;
      17'd11317: data = 8'he3;
      17'd11318: data = 8'he0;
      17'd11319: data = 8'he3;
      17'd11320: data = 8'he3;
      17'd11321: data = 8'he3;
      17'd11322: data = 8'he7;
      17'd11323: data = 8'he2;
      17'd11324: data = 8'hdb;
      17'd11325: data = 8'he2;
      17'd11326: data = 8'hde;
      17'd11327: data = 8'hd5;
      17'd11328: data = 8'hd3;
      17'd11329: data = 8'hd5;
      17'd11330: data = 8'hd3;
      17'd11331: data = 8'hcd;
      17'd11332: data = 8'hd2;
      17'd11333: data = 8'hd6;
      17'd11334: data = 8'hda;
      17'd11335: data = 8'hde;
      17'd11336: data = 8'he3;
      17'd11337: data = 8'hde;
      17'd11338: data = 8'hd3;
      17'd11339: data = 8'hd2;
      17'd11340: data = 8'hd2;
      17'd11341: data = 8'hd1;
      17'd11342: data = 8'hd5;
      17'd11343: data = 8'hdb;
      17'd11344: data = 8'he0;
      17'd11345: data = 8'hde;
      17'd11346: data = 8'he3;
      17'd11347: data = 8'heb;
      17'd11348: data = 8'he7;
      17'd11349: data = 8'he5;
      17'd11350: data = 8'he5;
      17'd11351: data = 8'he9;
      17'd11352: data = 8'he5;
      17'd11353: data = 8'he0;
      17'd11354: data = 8'heb;
      17'd11355: data = 8'hf4;
      17'd11356: data = 8'hf2;
      17'd11357: data = 8'hfa;
      17'd11358: data = 8'hfe;
      17'd11359: data = 8'hfe;
      17'd11360: data = 8'h00;
      17'd11361: data = 8'h01;
      17'd11362: data = 8'h01;
      17'd11363: data = 8'hfe;
      17'd11364: data = 8'h05;
      17'd11365: data = 8'h04;
      17'd11366: data = 8'h01;
      17'd11367: data = 8'h05;
      17'd11368: data = 8'h0a;
      17'd11369: data = 8'h0e;
      17'd11370: data = 8'h11;
      17'd11371: data = 8'h15;
      17'd11372: data = 8'h16;
      17'd11373: data = 8'h1b;
      17'd11374: data = 8'h16;
      17'd11375: data = 8'h13;
      17'd11376: data = 8'h19;
      17'd11377: data = 8'h11;
      17'd11378: data = 8'h13;
      17'd11379: data = 8'h13;
      17'd11380: data = 8'h12;
      17'd11381: data = 8'h1a;
      17'd11382: data = 8'h12;
      17'd11383: data = 8'h16;
      17'd11384: data = 8'h1e;
      17'd11385: data = 8'h1a;
      17'd11386: data = 8'h1e;
      17'd11387: data = 8'h15;
      17'd11388: data = 8'h12;
      17'd11389: data = 8'h11;
      17'd11390: data = 8'h0c;
      17'd11391: data = 8'h09;
      17'd11392: data = 8'h02;
      17'd11393: data = 8'h13;
      17'd11394: data = 8'h0c;
      17'd11395: data = 8'h02;
      17'd11396: data = 8'h1a;
      17'd11397: data = 8'h13;
      17'd11398: data = 8'h04;
      17'd11399: data = 8'h0a;
      17'd11400: data = 8'h00;
      17'd11401: data = 8'hfd;
      17'd11402: data = 8'hfe;
      17'd11403: data = 8'hfd;
      17'd11404: data = 8'hfe;
      17'd11405: data = 8'h01;
      17'd11406: data = 8'h0d;
      17'd11407: data = 8'hfd;
      17'd11408: data = 8'he5;
      17'd11409: data = 8'hf9;
      17'd11410: data = 8'h02;
      17'd11411: data = 8'h01;
      17'd11412: data = 8'h05;
      17'd11413: data = 8'h1a;
      17'd11414: data = 8'h1e;
      17'd11415: data = 8'hf4;
      17'd11416: data = 8'hda;
      17'd11417: data = 8'hdb;
      17'd11418: data = 8'hd3;
      17'd11419: data = 8'hc5;
      17'd11420: data = 8'he0;
      17'd11421: data = 8'h00;
      17'd11422: data = 8'h1a;
      17'd11423: data = 8'h23;
      17'd11424: data = 8'h23;
      17'd11425: data = 8'h23;
      17'd11426: data = 8'h12;
      17'd11427: data = 8'h02;
      17'd11428: data = 8'hf2;
      17'd11429: data = 8'hda;
      17'd11430: data = 8'hd1;
      17'd11431: data = 8'hd8;
      17'd11432: data = 8'hf2;
      17'd11433: data = 8'h05;
      17'd11434: data = 8'h13;
      17'd11435: data = 8'h43;
      17'd11436: data = 8'h52;
      17'd11437: data = 8'h2d;
      17'd11438: data = 8'h16;
      17'd11439: data = 8'h0a;
      17'd11440: data = 8'hf4;
      17'd11441: data = 8'hdb;
      17'd11442: data = 8'he9;
      17'd11443: data = 8'h0d;
      17'd11444: data = 8'h13;
      17'd11445: data = 8'h1b;
      17'd11446: data = 8'h2d;
      17'd11447: data = 8'h2f;
      17'd11448: data = 8'h24;
      17'd11449: data = 8'h22;
      17'd11450: data = 8'h26;
      17'd11451: data = 8'h0e;
      17'd11452: data = 8'h01;
      17'd11453: data = 8'h0c;
      17'd11454: data = 8'h09;
      17'd11455: data = 8'hfa;
      17'd11456: data = 8'h05;
      17'd11457: data = 8'h1c;
      17'd11458: data = 8'h1e;
      17'd11459: data = 8'h0d;
      17'd11460: data = 8'h0a;
      17'd11461: data = 8'h0d;
      17'd11462: data = 8'h0a;
      17'd11463: data = 8'hfc;
      17'd11464: data = 8'h05;
      17'd11465: data = 8'h13;
      17'd11466: data = 8'h01;
      17'd11467: data = 8'hf5;
      17'd11468: data = 8'hef;
      17'd11469: data = 8'he2;
      17'd11470: data = 8'hdb;
      17'd11471: data = 8'he3;
      17'd11472: data = 8'hed;
      17'd11473: data = 8'hef;
      17'd11474: data = 8'hfc;
      17'd11475: data = 8'h0a;
      17'd11476: data = 8'h00;
      17'd11477: data = 8'hef;
      17'd11478: data = 8'heb;
      17'd11479: data = 8'he9;
      17'd11480: data = 8'hdc;
      17'd11481: data = 8'hc9;
      17'd11482: data = 8'hce;
      17'd11483: data = 8'hda;
      17'd11484: data = 8'hde;
      17'd11485: data = 8'hf1;
      17'd11486: data = 8'h02;
      17'd11487: data = 8'h11;
      17'd11488: data = 8'h11;
      17'd11489: data = 8'h06;
      17'd11490: data = 8'hfc;
      17'd11491: data = 8'hed;
      17'd11492: data = 8'he4;
      17'd11493: data = 8'he5;
      17'd11494: data = 8'he7;
      17'd11495: data = 8'hf4;
      17'd11496: data = 8'h04;
      17'd11497: data = 8'h19;
      17'd11498: data = 8'h1f;
      17'd11499: data = 8'h1e;
      17'd11500: data = 8'h1f;
      17'd11501: data = 8'h23;
      17'd11502: data = 8'h1b;
      17'd11503: data = 8'h0c;
      17'd11504: data = 8'h0d;
      17'd11505: data = 8'h0e;
      17'd11506: data = 8'h0e;
      17'd11507: data = 8'h16;
      17'd11508: data = 8'h1a;
      17'd11509: data = 8'h26;
      17'd11510: data = 8'h2d;
      17'd11511: data = 8'h2b;
      17'd11512: data = 8'h29;
      17'd11513: data = 8'h27;
      17'd11514: data = 8'h24;
      17'd11515: data = 8'h22;
      17'd11516: data = 8'h1e;
      17'd11517: data = 8'h1e;
      17'd11518: data = 8'h23;
      17'd11519: data = 8'h27;
      17'd11520: data = 8'h22;
      17'd11521: data = 8'h16;
      17'd11522: data = 8'h12;
      17'd11523: data = 8'h13;
      17'd11524: data = 8'h12;
      17'd11525: data = 8'h0e;
      17'd11526: data = 8'h15;
      17'd11527: data = 8'h1e;
      17'd11528: data = 8'h1a;
      17'd11529: data = 8'h13;
      17'd11530: data = 8'h0e;
      17'd11531: data = 8'h06;
      17'd11532: data = 8'h00;
      17'd11533: data = 8'hf4;
      17'd11534: data = 8'hef;
      17'd11535: data = 8'hf2;
      17'd11536: data = 8'hf2;
      17'd11537: data = 8'hef;
      17'd11538: data = 8'hf1;
      17'd11539: data = 8'hf6;
      17'd11540: data = 8'hf5;
      17'd11541: data = 8'hf4;
      17'd11542: data = 8'heb;
      17'd11543: data = 8'hdc;
      17'd11544: data = 8'hdb;
      17'd11545: data = 8'hda;
      17'd11546: data = 8'hd8;
      17'd11547: data = 8'hd2;
      17'd11548: data = 8'hd8;
      17'd11549: data = 8'hde;
      17'd11550: data = 8'hda;
      17'd11551: data = 8'hd5;
      17'd11552: data = 8'hd2;
      17'd11553: data = 8'hd3;
      17'd11554: data = 8'hce;
      17'd11555: data = 8'hca;
      17'd11556: data = 8'hce;
      17'd11557: data = 8'hd2;
      17'd11558: data = 8'hcd;
      17'd11559: data = 8'hcd;
      17'd11560: data = 8'hd2;
      17'd11561: data = 8'hd5;
      17'd11562: data = 8'hd2;
      17'd11563: data = 8'hd3;
      17'd11564: data = 8'hd2;
      17'd11565: data = 8'hd3;
      17'd11566: data = 8'hd6;
      17'd11567: data = 8'hd5;
      17'd11568: data = 8'hda;
      17'd11569: data = 8'hdc;
      17'd11570: data = 8'he4;
      17'd11571: data = 8'he9;
      17'd11572: data = 8'he4;
      17'd11573: data = 8'he3;
      17'd11574: data = 8'he5;
      17'd11575: data = 8'he3;
      17'd11576: data = 8'hf4;
      17'd11577: data = 8'hf1;
      17'd11578: data = 8'hed;
      17'd11579: data = 8'h04;
      17'd11580: data = 8'hfa;
      17'd11581: data = 8'hf6;
      17'd11582: data = 8'h04;
      17'd11583: data = 8'hfe;
      17'd11584: data = 8'hf1;
      17'd11585: data = 8'hfc;
      17'd11586: data = 8'hf9;
      17'd11587: data = 8'hf9;
      17'd11588: data = 8'h0a;
      17'd11589: data = 8'h15;
      17'd11590: data = 8'h11;
      17'd11591: data = 8'h13;
      17'd11592: data = 8'h19;
      17'd11593: data = 8'h13;
      17'd11594: data = 8'h16;
      17'd11595: data = 8'h06;
      17'd11596: data = 8'h05;
      17'd11597: data = 8'h11;
      17'd11598: data = 8'h01;
      17'd11599: data = 8'h02;
      17'd11600: data = 8'h16;
      17'd11601: data = 8'h0d;
      17'd11602: data = 8'h0c;
      17'd11603: data = 8'h1b;
      17'd11604: data = 8'h13;
      17'd11605: data = 8'h16;
      17'd11606: data = 8'h24;
      17'd11607: data = 8'h19;
      17'd11608: data = 8'h12;
      17'd11609: data = 8'h16;
      17'd11610: data = 8'h13;
      17'd11611: data = 8'h0d;
      17'd11612: data = 8'h04;
      17'd11613: data = 8'h02;
      17'd11614: data = 8'h00;
      17'd11615: data = 8'hfc;
      17'd11616: data = 8'hf6;
      17'd11617: data = 8'h04;
      17'd11618: data = 8'h16;
      17'd11619: data = 8'h02;
      17'd11620: data = 8'h0c;
      17'd11621: data = 8'h23;
      17'd11622: data = 8'h05;
      17'd11623: data = 8'hfe;
      17'd11624: data = 8'h05;
      17'd11625: data = 8'hfd;
      17'd11626: data = 8'hfc;
      17'd11627: data = 8'hfc;
      17'd11628: data = 8'hfe;
      17'd11629: data = 8'hf4;
      17'd11630: data = 8'hfd;
      17'd11631: data = 8'h01;
      17'd11632: data = 8'hec;
      17'd11633: data = 8'hf4;
      17'd11634: data = 8'h05;
      17'd11635: data = 8'h02;
      17'd11636: data = 8'h0e;
      17'd11637: data = 8'h16;
      17'd11638: data = 8'h0d;
      17'd11639: data = 8'hf2;
      17'd11640: data = 8'he5;
      17'd11641: data = 8'he3;
      17'd11642: data = 8'hd3;
      17'd11643: data = 8'he2;
      17'd11644: data = 8'hf1;
      17'd11645: data = 8'hf4;
      17'd11646: data = 8'h09;
      17'd11647: data = 8'h19;
      17'd11648: data = 8'h19;
      17'd11649: data = 8'h1b;
      17'd11650: data = 8'h22;
      17'd11651: data = 8'h13;
      17'd11652: data = 8'h06;
      17'd11653: data = 8'h04;
      17'd11654: data = 8'he9;
      17'd11655: data = 8'he2;
      17'd11656: data = 8'hf4;
      17'd11657: data = 8'hfa;
      17'd11658: data = 8'h04;
      17'd11659: data = 8'h1f;
      17'd11660: data = 8'h29;
      17'd11661: data = 8'h1b;
      17'd11662: data = 8'h15;
      17'd11663: data = 8'h23;
      17'd11664: data = 8'h11;
      17'd11665: data = 8'h0a;
      17'd11666: data = 8'h24;
      17'd11667: data = 8'h1e;
      17'd11668: data = 8'h0c;
      17'd11669: data = 8'h0e;
      17'd11670: data = 8'h0c;
      17'd11671: data = 8'hfc;
      17'd11672: data = 8'h04;
      17'd11673: data = 8'h16;
      17'd11674: data = 8'h11;
      17'd11675: data = 8'h19;
      17'd11676: data = 8'h19;
      17'd11677: data = 8'h16;
      17'd11678: data = 8'h1c;
      17'd11679: data = 8'h16;
      17'd11680: data = 8'h16;
      17'd11681: data = 8'h19;
      17'd11682: data = 8'h0a;
      17'd11683: data = 8'hf6;
      17'd11684: data = 8'heb;
      17'd11685: data = 8'heb;
      17'd11686: data = 8'he5;
      17'd11687: data = 8'he9;
      17'd11688: data = 8'hfe;
      17'd11689: data = 8'h01;
      17'd11690: data = 8'h00;
      17'd11691: data = 8'hfe;
      17'd11692: data = 8'hf6;
      17'd11693: data = 8'hed;
      17'd11694: data = 8'he3;
      17'd11695: data = 8'he7;
      17'd11696: data = 8'hde;
      17'd11697: data = 8'hd8;
      17'd11698: data = 8'hde;
      17'd11699: data = 8'hdc;
      17'd11700: data = 8'hdb;
      17'd11701: data = 8'he0;
      17'd11702: data = 8'he5;
      17'd11703: data = 8'heb;
      17'd11704: data = 8'he9;
      17'd11705: data = 8'he9;
      17'd11706: data = 8'heb;
      17'd11707: data = 8'he7;
      17'd11708: data = 8'hed;
      17'd11709: data = 8'hf1;
      17'd11710: data = 8'hf4;
      17'd11711: data = 8'hfd;
      17'd11712: data = 8'hfd;
      17'd11713: data = 8'hf6;
      17'd11714: data = 8'hfa;
      17'd11715: data = 8'hf9;
      17'd11716: data = 8'hf6;
      17'd11717: data = 8'h02;
      17'd11718: data = 8'h0c;
      17'd11719: data = 8'h0d;
      17'd11720: data = 8'h1b;
      17'd11721: data = 8'h26;
      17'd11722: data = 8'h27;
      17'd11723: data = 8'h27;
      17'd11724: data = 8'h27;
      17'd11725: data = 8'h23;
      17'd11726: data = 8'h1b;
      17'd11727: data = 8'h1a;
      17'd11728: data = 8'h1b;
      17'd11729: data = 8'h1c;
      17'd11730: data = 8'h26;
      17'd11731: data = 8'h2d;
      17'd11732: data = 8'h33;
      17'd11733: data = 8'h39;
      17'd11734: data = 8'h39;
      17'd11735: data = 8'h34;
      17'd11736: data = 8'h2f;
      17'd11737: data = 8'h2d;
      17'd11738: data = 8'h29;
      17'd11739: data = 8'h24;
      17'd11740: data = 8'h27;
      17'd11741: data = 8'h24;
      17'd11742: data = 8'h26;
      17'd11743: data = 8'h2b;
      17'd11744: data = 8'h1f;
      17'd11745: data = 8'h1a;
      17'd11746: data = 8'h19;
      17'd11747: data = 8'h11;
      17'd11748: data = 8'h0c;
      17'd11749: data = 8'h12;
      17'd11750: data = 8'h0e;
      17'd11751: data = 8'h06;
      17'd11752: data = 8'h0c;
      17'd11753: data = 8'h09;
      17'd11754: data = 8'h02;
      17'd11755: data = 8'h02;
      17'd11756: data = 8'h00;
      17'd11757: data = 8'hf4;
      17'd11758: data = 8'hec;
      17'd11759: data = 8'he7;
      17'd11760: data = 8'he3;
      17'd11761: data = 8'hde;
      17'd11762: data = 8'he2;
      17'd11763: data = 8'he2;
      17'd11764: data = 8'hdc;
      17'd11765: data = 8'hde;
      17'd11766: data = 8'hda;
      17'd11767: data = 8'hd8;
      17'd11768: data = 8'hd3;
      17'd11769: data = 8'hd1;
      17'd11770: data = 8'hce;
      17'd11771: data = 8'hce;
      17'd11772: data = 8'hd1;
      17'd11773: data = 8'hcd;
      17'd11774: data = 8'hcd;
      17'd11775: data = 8'hd1;
      17'd11776: data = 8'hca;
      17'd11777: data = 8'hca;
      17'd11778: data = 8'hcb;
      17'd11779: data = 8'hc4;
      17'd11780: data = 8'hc4;
      17'd11781: data = 8'hc6;
      17'd11782: data = 8'hcd;
      17'd11783: data = 8'hce;
      17'd11784: data = 8'hd6;
      17'd11785: data = 8'he0;
      17'd11786: data = 8'hdb;
      17'd11787: data = 8'hde;
      17'd11788: data = 8'hdc;
      17'd11789: data = 8'hd6;
      17'd11790: data = 8'hda;
      17'd11791: data = 8'hdc;
      17'd11792: data = 8'he3;
      17'd11793: data = 8'he7;
      17'd11794: data = 8'heb;
      17'd11795: data = 8'hed;
      17'd11796: data = 8'hf1;
      17'd11797: data = 8'hf5;
      17'd11798: data = 8'hf5;
      17'd11799: data = 8'hf2;
      17'd11800: data = 8'hf9;
      17'd11801: data = 8'hfa;
      17'd11802: data = 8'hfd;
      17'd11803: data = 8'h04;
      17'd11804: data = 8'h06;
      17'd11805: data = 8'h09;
      17'd11806: data = 8'h09;
      17'd11807: data = 8'h0a;
      17'd11808: data = 8'h04;
      17'd11809: data = 8'h04;
      17'd11810: data = 8'h05;
      17'd11811: data = 8'h02;
      17'd11812: data = 8'h06;
      17'd11813: data = 8'h09;
      17'd11814: data = 8'h0c;
      17'd11815: data = 8'h12;
      17'd11816: data = 8'h19;
      17'd11817: data = 8'h1a;
      17'd11818: data = 8'h15;
      17'd11819: data = 8'h12;
      17'd11820: data = 8'h0c;
      17'd11821: data = 8'h05;
      17'd11822: data = 8'h0a;
      17'd11823: data = 8'h0a;
      17'd11824: data = 8'h09;
      17'd11825: data = 8'h12;
      17'd11826: data = 8'h0d;
      17'd11827: data = 8'h0a;
      17'd11828: data = 8'h09;
      17'd11829: data = 8'h06;
      17'd11830: data = 8'h05;
      17'd11831: data = 8'h01;
      17'd11832: data = 8'h04;
      17'd11833: data = 8'h05;
      17'd11834: data = 8'h05;
      17'd11835: data = 8'h06;
      17'd11836: data = 8'h02;
      17'd11837: data = 8'h02;
      17'd11838: data = 8'h04;
      17'd11839: data = 8'h00;
      17'd11840: data = 8'h01;
      17'd11841: data = 8'h04;
      17'd11842: data = 8'hfa;
      17'd11843: data = 8'hef;
      17'd11844: data = 8'hfe;
      17'd11845: data = 8'h06;
      17'd11846: data = 8'hf9;
      17'd11847: data = 8'h01;
      17'd11848: data = 8'h09;
      17'd11849: data = 8'h02;
      17'd11850: data = 8'hfd;
      17'd11851: data = 8'hf4;
      17'd11852: data = 8'h00;
      17'd11853: data = 8'h0c;
      17'd11854: data = 8'hfd;
      17'd11855: data = 8'h00;
      17'd11856: data = 8'h06;
      17'd11857: data = 8'hfe;
      17'd11858: data = 8'hfd;
      17'd11859: data = 8'h02;
      17'd11860: data = 8'hfc;
      17'd11861: data = 8'hfa;
      17'd11862: data = 8'h0a;
      17'd11863: data = 8'h09;
      17'd11864: data = 8'he4;
      17'd11865: data = 8'hd5;
      17'd11866: data = 8'hf4;
      17'd11867: data = 8'h06;
      17'd11868: data = 8'hf4;
      17'd11869: data = 8'h06;
      17'd11870: data = 8'h3a;
      17'd11871: data = 8'h2b;
      17'd11872: data = 8'h0c;
      17'd11873: data = 8'h16;
      17'd11874: data = 8'h1a;
      17'd11875: data = 8'h0c;
      17'd11876: data = 8'h02;
      17'd11877: data = 8'h06;
      17'd11878: data = 8'h11;
      17'd11879: data = 8'h04;
      17'd11880: data = 8'h01;
      17'd11881: data = 8'h09;
      17'd11882: data = 8'h01;
      17'd11883: data = 8'h09;
      17'd11884: data = 8'h2c;
      17'd11885: data = 8'h26;
      17'd11886: data = 8'h00;
      17'd11887: data = 8'h0a;
      17'd11888: data = 8'h27;
      17'd11889: data = 8'h1b;
      17'd11890: data = 8'h09;
      17'd11891: data = 8'h1f;
      17'd11892: data = 8'h43;
      17'd11893: data = 8'h22;
      17'd11894: data = 8'hf6;
      17'd11895: data = 8'h0c;
      17'd11896: data = 8'h0a;
      17'd11897: data = 8'hf2;
      17'd11898: data = 8'hfd;
      17'd11899: data = 8'h0e;
      17'd11900: data = 8'h0d;
      17'd11901: data = 8'h0a;
      17'd11902: data = 8'h0c;
      17'd11903: data = 8'h02;
      17'd11904: data = 8'hf6;
      17'd11905: data = 8'h01;
      17'd11906: data = 8'h15;
      17'd11907: data = 8'hfd;
      17'd11908: data = 8'hde;
      17'd11909: data = 8'hf4;
      17'd11910: data = 8'hfc;
      17'd11911: data = 8'hdc;
      17'd11912: data = 8'hd6;
      17'd11913: data = 8'hf1;
      17'd11914: data = 8'hfa;
      17'd11915: data = 8'he2;
      17'd11916: data = 8'hcb;
      17'd11917: data = 8'hd8;
      17'd11918: data = 8'hdb;
      17'd11919: data = 8'hca;
      17'd11920: data = 8'hd3;
      17'd11921: data = 8'hec;
      17'd11922: data = 8'hed;
      17'd11923: data = 8'hf4;
      17'd11924: data = 8'hf4;
      17'd11925: data = 8'he3;
      17'd11926: data = 8'he0;
      17'd11927: data = 8'hed;
      17'd11928: data = 8'hef;
      17'd11929: data = 8'he5;
      17'd11930: data = 8'he0;
      17'd11931: data = 8'hf5;
      17'd11932: data = 8'h01;
      17'd11933: data = 8'hf1;
      17'd11934: data = 8'hf5;
      17'd11935: data = 8'h0e;
      17'd11936: data = 8'h13;
      17'd11937: data = 8'h06;
      17'd11938: data = 8'h05;
      17'd11939: data = 8'h13;
      17'd11940: data = 8'h1f;
      17'd11941: data = 8'h19;
      17'd11942: data = 8'h1b;
      17'd11943: data = 8'h2f;
      17'd11944: data = 8'h35;
      17'd11945: data = 8'h31;
      17'd11946: data = 8'h31;
      17'd11947: data = 8'h27;
      17'd11948: data = 8'h27;
      17'd11949: data = 8'h2c;
      17'd11950: data = 8'h27;
      17'd11951: data = 8'h23;
      17'd11952: data = 8'h29;
      17'd11953: data = 8'h35;
      17'd11954: data = 8'h3d;
      17'd11955: data = 8'h34;
      17'd11956: data = 8'h2d;
      17'd11957: data = 8'h3e;
      17'd11958: data = 8'h3d;
      17'd11959: data = 8'h2c;
      17'd11960: data = 8'h27;
      17'd11961: data = 8'h31;
      17'd11962: data = 8'h2f;
      17'd11963: data = 8'h23;
      17'd11964: data = 8'h1c;
      17'd11965: data = 8'h29;
      17'd11966: data = 8'h27;
      17'd11967: data = 8'h12;
      17'd11968: data = 8'h0e;
      17'd11969: data = 8'h0a;
      17'd11970: data = 8'h00;
      17'd11971: data = 8'h04;
      17'd11972: data = 8'h05;
      17'd11973: data = 8'hfe;
      17'd11974: data = 8'h02;
      17'd11975: data = 8'h0c;
      17'd11976: data = 8'h04;
      17'd11977: data = 8'hf5;
      17'd11978: data = 8'hef;
      17'd11979: data = 8'hf4;
      17'd11980: data = 8'hec;
      17'd11981: data = 8'hd6;
      17'd11982: data = 8'hd6;
      17'd11983: data = 8'he3;
      17'd11984: data = 8'hd8;
      17'd11985: data = 8'hce;
      17'd11986: data = 8'hd5;
      17'd11987: data = 8'hda;
      17'd11988: data = 8'hd5;
      17'd11989: data = 8'hcd;
      17'd11990: data = 8'hce;
      17'd11991: data = 8'hd2;
      17'd11992: data = 8'hc9;
      17'd11993: data = 8'hcd;
      17'd11994: data = 8'hd3;
      17'd11995: data = 8'hd1;
      17'd11996: data = 8'hd6;
      17'd11997: data = 8'hdc;
      17'd11998: data = 8'hd2;
      17'd11999: data = 8'hca;
      17'd12000: data = 8'hce;
      17'd12001: data = 8'hd3;
      17'd12002: data = 8'hc9;
      17'd12003: data = 8'hc5;
      17'd12004: data = 8'hd3;
      17'd12005: data = 8'hde;
      17'd12006: data = 8'hd8;
      17'd12007: data = 8'hda;
      17'd12008: data = 8'he7;
      17'd12009: data = 8'he7;
      17'd12010: data = 8'he5;
      17'd12011: data = 8'he9;
      17'd12012: data = 8'heb;
      17'd12013: data = 8'hed;
      17'd12014: data = 8'hf2;
      17'd12015: data = 8'hf9;
      17'd12016: data = 8'hfe;
      17'd12017: data = 8'hfc;
      17'd12018: data = 8'hfc;
      17'd12019: data = 8'h01;
      17'd12020: data = 8'hf9;
      17'd12021: data = 8'hf4;
      17'd12022: data = 8'hfc;
      17'd12023: data = 8'hfe;
      17'd12024: data = 8'hfd;
      17'd12025: data = 8'h01;
      17'd12026: data = 8'h09;
      17'd12027: data = 8'h0e;
      17'd12028: data = 8'h0c;
      17'd12029: data = 8'h0a;
      17'd12030: data = 8'h0e;
      17'd12031: data = 8'h0a;
      17'd12032: data = 8'h00;
      17'd12033: data = 8'h02;
      17'd12034: data = 8'h05;
      17'd12035: data = 8'h04;
      17'd12036: data = 8'h0a;
      17'd12037: data = 8'h0c;
      17'd12038: data = 8'h0a;
      17'd12039: data = 8'h09;
      17'd12040: data = 8'h09;
      17'd12041: data = 8'h05;
      17'd12042: data = 8'h00;
      17'd12043: data = 8'hfd;
      17'd12044: data = 8'h01;
      17'd12045: data = 8'h05;
      17'd12046: data = 8'h01;
      17'd12047: data = 8'h06;
      17'd12048: data = 8'h0d;
      17'd12049: data = 8'h06;
      17'd12050: data = 8'h04;
      17'd12051: data = 8'h02;
      17'd12052: data = 8'h02;
      17'd12053: data = 8'hfc;
      17'd12054: data = 8'hf4;
      17'd12055: data = 8'hfa;
      17'd12056: data = 8'hfe;
      17'd12057: data = 8'h00;
      17'd12058: data = 8'h01;
      17'd12059: data = 8'h01;
      17'd12060: data = 8'h02;
      17'd12061: data = 8'h01;
      17'd12062: data = 8'hf6;
      17'd12063: data = 8'hfe;
      17'd12064: data = 8'hfe;
      17'd12065: data = 8'hfa;
      17'd12066: data = 8'hfe;
      17'd12067: data = 8'h04;
      17'd12068: data = 8'h01;
      17'd12069: data = 8'h01;
      17'd12070: data = 8'h05;
      17'd12071: data = 8'h02;
      17'd12072: data = 8'h01;
      17'd12073: data = 8'h02;
      17'd12074: data = 8'h02;
      17'd12075: data = 8'h01;
      17'd12076: data = 8'h01;
      17'd12077: data = 8'h02;
      17'd12078: data = 8'h0d;
      17'd12079: data = 8'h12;
      17'd12080: data = 8'h11;
      17'd12081: data = 8'h13;
      17'd12082: data = 8'hfd;
      17'd12083: data = 8'he4;
      17'd12084: data = 8'hde;
      17'd12085: data = 8'hde;
      17'd12086: data = 8'he0;
      17'd12087: data = 8'hf1;
      17'd12088: data = 8'hfe;
      17'd12089: data = 8'h16;
      17'd12090: data = 8'h1c;
      17'd12091: data = 8'h0e;
      17'd12092: data = 8'h0d;
      17'd12093: data = 8'h0e;
      17'd12094: data = 8'h06;
      17'd12095: data = 8'h12;
      17'd12096: data = 8'h1e;
      17'd12097: data = 8'h1a;
      17'd12098: data = 8'h1a;
      17'd12099: data = 8'h0e;
      17'd12100: data = 8'h0c;
      17'd12101: data = 8'h12;
      17'd12102: data = 8'h0c;
      17'd12103: data = 8'h0c;
      17'd12104: data = 8'h06;
      17'd12105: data = 8'hfa;
      17'd12106: data = 8'hf9;
      17'd12107: data = 8'hfe;
      17'd12108: data = 8'hfd;
      17'd12109: data = 8'h0d;
      17'd12110: data = 8'h29;
      17'd12111: data = 8'h34;
      17'd12112: data = 8'h34;
      17'd12113: data = 8'h23;
      17'd12114: data = 8'h12;
      17'd12115: data = 8'h11;
      17'd12116: data = 8'h02;
      17'd12117: data = 8'h0a;
      17'd12118: data = 8'h22;
      17'd12119: data = 8'h1f;
      17'd12120: data = 8'h13;
      17'd12121: data = 8'h0a;
      17'd12122: data = 8'hfe;
      17'd12123: data = 8'hf6;
      17'd12124: data = 8'hf1;
      17'd12125: data = 8'heb;
      17'd12126: data = 8'hf2;
      17'd12127: data = 8'hef;
      17'd12128: data = 8'he9;
      17'd12129: data = 8'hed;
      17'd12130: data = 8'hec;
      17'd12131: data = 8'hf1;
      17'd12132: data = 8'h00;
      17'd12133: data = 8'h01;
      17'd12134: data = 8'hf9;
      17'd12135: data = 8'hed;
      17'd12136: data = 8'hdb;
      17'd12137: data = 8'hce;
      17'd12138: data = 8'hca;
      17'd12139: data = 8'hcb;
      17'd12140: data = 8'he0;
      17'd12141: data = 8'he4;
      17'd12142: data = 8'hdb;
      17'd12143: data = 8'hda;
      17'd12144: data = 8'hd1;
      17'd12145: data = 8'hca;
      17'd12146: data = 8'hce;
      17'd12147: data = 8'hd3;
      17'd12148: data = 8'he3;
      17'd12149: data = 8'hf1;
      17'd12150: data = 8'hf1;
      17'd12151: data = 8'hf6;
      17'd12152: data = 8'hfa;
      17'd12153: data = 8'hfe;
      17'd12154: data = 8'h0a;
      17'd12155: data = 8'h0c;
      17'd12156: data = 8'h0c;
      17'd12157: data = 8'h0a;
      17'd12158: data = 8'h01;
      17'd12159: data = 8'hfe;
      17'd12160: data = 8'h01;
      17'd12161: data = 8'h0c;
      17'd12162: data = 8'h22;
      17'd12163: data = 8'h2b;
      17'd12164: data = 8'h29;
      17'd12165: data = 8'h2c;
      17'd12166: data = 8'h29;
      17'd12167: data = 8'h23;
      17'd12168: data = 8'h26;
      17'd12169: data = 8'h2c;
      17'd12170: data = 8'h36;
      17'd12171: data = 8'h3e;
      17'd12172: data = 8'h40;
      17'd12173: data = 8'h43;
      17'd12174: data = 8'h3e;
      17'd12175: data = 8'h36;
      17'd12176: data = 8'h35;
      17'd12177: data = 8'h39;
      17'd12178: data = 8'h34;
      17'd12179: data = 8'h31;
      17'd12180: data = 8'h2c;
      17'd12181: data = 8'h24;
      17'd12182: data = 8'h24;
      17'd12183: data = 8'h24;
      17'd12184: data = 8'h29;
      17'd12185: data = 8'h2b;
      17'd12186: data = 8'h22;
      17'd12187: data = 8'h1c;
      17'd12188: data = 8'h16;
      17'd12189: data = 8'h09;
      17'd12190: data = 8'h09;
      17'd12191: data = 8'h0d;
      17'd12192: data = 8'h0e;
      17'd12193: data = 8'h12;
      17'd12194: data = 8'h0d;
      17'd12195: data = 8'h09;
      17'd12196: data = 8'h00;
      17'd12197: data = 8'hf2;
      17'd12198: data = 8'hef;
      17'd12199: data = 8'hed;
      17'd12200: data = 8'he7;
      17'd12201: data = 8'he7;
      17'd12202: data = 8'he7;
      17'd12203: data = 8'hdc;
      17'd12204: data = 8'hda;
      17'd12205: data = 8'hd8;
      17'd12206: data = 8'hd5;
      17'd12207: data = 8'hd5;
      17'd12208: data = 8'hd3;
      17'd12209: data = 8'hce;
      17'd12210: data = 8'hce;
      17'd12211: data = 8'hca;
      17'd12212: data = 8'hce;
      17'd12213: data = 8'hd8;
      17'd12214: data = 8'hd8;
      17'd12215: data = 8'hdc;
      17'd12216: data = 8'hde;
      17'd12217: data = 8'hd8;
      17'd12218: data = 8'hd2;
      17'd12219: data = 8'hce;
      17'd12220: data = 8'hce;
      17'd12221: data = 8'hd5;
      17'd12222: data = 8'hd6;
      17'd12223: data = 8'hdb;
      17'd12224: data = 8'he0;
      17'd12225: data = 8'hde;
      17'd12226: data = 8'hdc;
      17'd12227: data = 8'hdc;
      17'd12228: data = 8'hdc;
      17'd12229: data = 8'he2;
      17'd12230: data = 8'he7;
      17'd12231: data = 8'he9;
      17'd12232: data = 8'hf1;
      17'd12233: data = 8'hf2;
      17'd12234: data = 8'hf6;
      17'd12235: data = 8'hfd;
      17'd12236: data = 8'hfe;
      17'd12237: data = 8'h02;
      17'd12238: data = 8'h01;
      17'd12239: data = 8'hfd;
      17'd12240: data = 8'hfd;
      17'd12241: data = 8'h00;
      17'd12242: data = 8'h02;
      17'd12243: data = 8'h09;
      17'd12244: data = 8'h0c;
      17'd12245: data = 8'h0c;
      17'd12246: data = 8'h09;
      17'd12247: data = 8'h06;
      17'd12248: data = 8'h04;
      17'd12249: data = 8'h01;
      17'd12250: data = 8'h04;
      17'd12251: data = 8'h04;
      17'd12252: data = 8'h05;
      17'd12253: data = 8'h05;
      17'd12254: data = 8'h06;
      17'd12255: data = 8'h09;
      17'd12256: data = 8'h09;
      17'd12257: data = 8'h0a;
      17'd12258: data = 8'h09;
      17'd12259: data = 8'h05;
      17'd12260: data = 8'h02;
      17'd12261: data = 8'hfd;
      17'd12262: data = 8'hfd;
      17'd12263: data = 8'hfe;
      17'd12264: data = 8'hfd;
      17'd12265: data = 8'h00;
      17'd12266: data = 8'h00;
      17'd12267: data = 8'h01;
      17'd12268: data = 8'hfe;
      17'd12269: data = 8'hfc;
      17'd12270: data = 8'hf9;
      17'd12271: data = 8'hfa;
      17'd12272: data = 8'hfc;
      17'd12273: data = 8'hfa;
      17'd12274: data = 8'hfa;
      17'd12275: data = 8'hfa;
      17'd12276: data = 8'hf9;
      17'd12277: data = 8'hfc;
      17'd12278: data = 8'h00;
      17'd12279: data = 8'hfd;
      17'd12280: data = 8'h00;
      17'd12281: data = 8'hf9;
      17'd12282: data = 8'hfc;
      17'd12283: data = 8'hf9;
      17'd12284: data = 8'hf4;
      17'd12285: data = 8'h00;
      17'd12286: data = 8'h02;
      17'd12287: data = 8'h00;
      17'd12288: data = 8'hfe;
      17'd12289: data = 8'h04;
      17'd12290: data = 8'hfe;
      17'd12291: data = 8'hfd;
      17'd12292: data = 8'h02;
      17'd12293: data = 8'h02;
      17'd12294: data = 8'h05;
      17'd12295: data = 8'h05;
      17'd12296: data = 8'h06;
      17'd12297: data = 8'h0c;
      17'd12298: data = 8'h04;
      17'd12299: data = 8'h09;
      17'd12300: data = 8'h11;
      17'd12301: data = 8'h0e;
      17'd12302: data = 8'h0e;
      17'd12303: data = 8'h15;
      17'd12304: data = 8'h15;
      17'd12305: data = 8'h05;
      17'd12306: data = 8'hf6;
      17'd12307: data = 8'hf4;
      17'd12308: data = 8'h01;
      17'd12309: data = 8'hf5;
      17'd12310: data = 8'heb;
      17'd12311: data = 8'hfc;
      17'd12312: data = 8'h01;
      17'd12313: data = 8'hf9;
      17'd12314: data = 8'hf4;
      17'd12315: data = 8'h02;
      17'd12316: data = 8'h00;
      17'd12317: data = 8'hf9;
      17'd12318: data = 8'h02;
      17'd12319: data = 8'h15;
      17'd12320: data = 8'h15;
      17'd12321: data = 8'h09;
      17'd12322: data = 8'h1a;
      17'd12323: data = 8'h16;
      17'd12324: data = 8'h0c;
      17'd12325: data = 8'h15;
      17'd12326: data = 8'h1e;
      17'd12327: data = 8'h0e;
      17'd12328: data = 8'hfd;
      17'd12329: data = 8'h06;
      17'd12330: data = 8'h0e;
      17'd12331: data = 8'h01;
      17'd12332: data = 8'hfc;
      17'd12333: data = 8'h0e;
      17'd12334: data = 8'h12;
      17'd12335: data = 8'h01;
      17'd12336: data = 8'h02;
      17'd12337: data = 8'h0a;
      17'd12338: data = 8'h05;
      17'd12339: data = 8'h01;
      17'd12340: data = 8'h11;
      17'd12341: data = 8'h1f;
      17'd12342: data = 8'h16;
      17'd12343: data = 8'h12;
      17'd12344: data = 8'h1a;
      17'd12345: data = 8'h11;
      17'd12346: data = 8'h04;
      17'd12347: data = 8'h06;
      17'd12348: data = 8'h0d;
      17'd12349: data = 8'h00;
      17'd12350: data = 8'hf4;
      17'd12351: data = 8'hfa;
      17'd12352: data = 8'hf6;
      17'd12353: data = 8'he3;
      17'd12354: data = 8'he3;
      17'd12355: data = 8'hf2;
      17'd12356: data = 8'he9;
      17'd12357: data = 8'hdc;
      17'd12358: data = 8'hdb;
      17'd12359: data = 8'he2;
      17'd12360: data = 8'hd6;
      17'd12361: data = 8'hd1;
      17'd12362: data = 8'he4;
      17'd12363: data = 8'hed;
      17'd12364: data = 8'he9;
      17'd12365: data = 8'he7;
      17'd12366: data = 8'he9;
      17'd12367: data = 8'he4;
      17'd12368: data = 8'he2;
      17'd12369: data = 8'he5;
      17'd12370: data = 8'he7;
      17'd12371: data = 8'he5;
      17'd12372: data = 8'he2;
      17'd12373: data = 8'he7;
      17'd12374: data = 8'heb;
      17'd12375: data = 8'he4;
      17'd12376: data = 8'heb;
      17'd12377: data = 8'hf4;
      17'd12378: data = 8'hf9;
      17'd12379: data = 8'hf9;
      17'd12380: data = 8'hf6;
      17'd12381: data = 8'hfe;
      17'd12382: data = 8'h04;
      17'd12383: data = 8'h04;
      17'd12384: data = 8'h0d;
      17'd12385: data = 8'h23;
      17'd12386: data = 8'h26;
      17'd12387: data = 8'h23;
      17'd12388: data = 8'h27;
      17'd12389: data = 8'h29;
      17'd12390: data = 8'h24;
      17'd12391: data = 8'h26;
      17'd12392: data = 8'h2c;
      17'd12393: data = 8'h33;
      17'd12394: data = 8'h2b;
      17'd12395: data = 8'h2d;
      17'd12396: data = 8'h2f;
      17'd12397: data = 8'h29;
      17'd12398: data = 8'h26;
      17'd12399: data = 8'h2d;
      17'd12400: data = 8'h2d;
      17'd12401: data = 8'h27;
      17'd12402: data = 8'h26;
      17'd12403: data = 8'h29;
      17'd12404: data = 8'h2b;
      17'd12405: data = 8'h1f;
      17'd12406: data = 8'h26;
      17'd12407: data = 8'h33;
      17'd12408: data = 8'h2c;
      17'd12409: data = 8'h26;
      17'd12410: data = 8'h27;
      17'd12411: data = 8'h26;
      17'd12412: data = 8'h19;
      17'd12413: data = 8'h16;
      17'd12414: data = 8'h16;
      17'd12415: data = 8'h12;
      17'd12416: data = 8'h0c;
      17'd12417: data = 8'h06;
      17'd12418: data = 8'h0c;
      17'd12419: data = 8'hfd;
      17'd12420: data = 8'hef;
      17'd12421: data = 8'hf4;
      17'd12422: data = 8'hf2;
      17'd12423: data = 8'he5;
      17'd12424: data = 8'he4;
      17'd12425: data = 8'heb;
      17'd12426: data = 8'he5;
      17'd12427: data = 8'he0;
      17'd12428: data = 8'he3;
      17'd12429: data = 8'heb;
      17'd12430: data = 8'he4;
      17'd12431: data = 8'hda;
      17'd12432: data = 8'hdc;
      17'd12433: data = 8'hda;
      17'd12434: data = 8'hd1;
      17'd12435: data = 8'hd3;
      17'd12436: data = 8'hd8;
      17'd12437: data = 8'hd5;
      17'd12438: data = 8'hd3;
      17'd12439: data = 8'hdb;
      17'd12440: data = 8'hda;
      17'd12441: data = 8'hd1;
      17'd12442: data = 8'hcd;
      17'd12443: data = 8'hd3;
      17'd12444: data = 8'hd5;
      17'd12445: data = 8'hce;
      17'd12446: data = 8'hd6;
      17'd12447: data = 8'hde;
      17'd12448: data = 8'hdc;
      17'd12449: data = 8'he0;
      17'd12450: data = 8'he4;
      17'd12451: data = 8'heb;
      17'd12452: data = 8'he9;
      17'd12453: data = 8'heb;
      17'd12454: data = 8'hed;
      17'd12455: data = 8'hed;
      17'd12456: data = 8'hed;
      17'd12457: data = 8'hf4;
      17'd12458: data = 8'hfc;
      17'd12459: data = 8'hf9;
      17'd12460: data = 8'hfd;
      17'd12461: data = 8'h01;
      17'd12462: data = 8'hfe;
      17'd12463: data = 8'hfc;
      17'd12464: data = 8'h00;
      17'd12465: data = 8'h06;
      17'd12466: data = 8'h05;
      17'd12467: data = 8'h04;
      17'd12468: data = 8'h04;
      17'd12469: data = 8'h0a;
      17'd12470: data = 8'h0a;
      17'd12471: data = 8'h09;
      17'd12472: data = 8'h0d;
      17'd12473: data = 8'h0c;
      17'd12474: data = 8'h0a;
      17'd12475: data = 8'h06;
      17'd12476: data = 8'h06;
      17'd12477: data = 8'h09;
      17'd12478: data = 8'h05;
      17'd12479: data = 8'h09;
      17'd12480: data = 8'h0a;
      17'd12481: data = 8'h04;
      17'd12482: data = 8'h00;
      17'd12483: data = 8'h00;
      17'd12484: data = 8'hfd;
      17'd12485: data = 8'hf5;
      17'd12486: data = 8'hfa;
      17'd12487: data = 8'h00;
      17'd12488: data = 8'hfc;
      17'd12489: data = 8'hfa;
      17'd12490: data = 8'hfd;
      17'd12491: data = 8'hfe;
      17'd12492: data = 8'hf9;
      17'd12493: data = 8'hf9;
      17'd12494: data = 8'hfc;
      17'd12495: data = 8'hfc;
      17'd12496: data = 8'hfa;
      17'd12497: data = 8'hfa;
      17'd12498: data = 8'hfd;
      17'd12499: data = 8'hf6;
      17'd12500: data = 8'hfa;
      17'd12501: data = 8'hfe;
      17'd12502: data = 8'h01;
      17'd12503: data = 8'hfd;
      17'd12504: data = 8'hf9;
      17'd12505: data = 8'hf6;
      17'd12506: data = 8'hf9;
      17'd12507: data = 8'hf6;
      17'd12508: data = 8'hfe;
      17'd12509: data = 8'h00;
      17'd12510: data = 8'hfd;
      17'd12511: data = 8'h0a;
      17'd12512: data = 8'hfd;
      17'd12513: data = 8'h02;
      17'd12514: data = 8'h04;
      17'd12515: data = 8'h01;
      17'd12516: data = 8'h04;
      17'd12517: data = 8'h00;
      17'd12518: data = 8'h0d;
      17'd12519: data = 8'h06;
      17'd12520: data = 8'h04;
      17'd12521: data = 8'h0e;
      17'd12522: data = 8'h0c;
      17'd12523: data = 8'h0e;
      17'd12524: data = 8'h0e;
      17'd12525: data = 8'h12;
      17'd12526: data = 8'h0d;
      17'd12527: data = 8'h0a;
      17'd12528: data = 8'h0d;
      17'd12529: data = 8'h12;
      17'd12530: data = 8'h0d;
      17'd12531: data = 8'h11;
      17'd12532: data = 8'h0e;
      17'd12533: data = 8'hfe;
      17'd12534: data = 8'h01;
      17'd12535: data = 8'hfa;
      17'd12536: data = 8'hf6;
      17'd12537: data = 8'hf6;
      17'd12538: data = 8'hf2;
      17'd12539: data = 8'hfe;
      17'd12540: data = 8'hf6;
      17'd12541: data = 8'hf4;
      17'd12542: data = 8'hf4;
      17'd12543: data = 8'hfa;
      17'd12544: data = 8'h01;
      17'd12545: data = 8'hfe;
      17'd12546: data = 8'h06;
      17'd12547: data = 8'h04;
      17'd12548: data = 8'h09;
      17'd12549: data = 8'h0a;
      17'd12550: data = 8'h0a;
      17'd12551: data = 8'h12;
      17'd12552: data = 8'h19;
      17'd12553: data = 8'h1a;
      17'd12554: data = 8'h15;
      17'd12555: data = 8'h0c;
      17'd12556: data = 8'h06;
      17'd12557: data = 8'h06;
      17'd12558: data = 8'h01;
      17'd12559: data = 8'h04;
      17'd12560: data = 8'h0d;
      17'd12561: data = 8'h05;
      17'd12562: data = 8'h09;
      17'd12563: data = 8'h04;
      17'd12564: data = 8'h00;
      17'd12565: data = 8'h06;
      17'd12566: data = 8'h04;
      17'd12567: data = 8'h06;
      17'd12568: data = 8'h09;
      17'd12569: data = 8'h09;
      17'd12570: data = 8'h0d;
      17'd12571: data = 8'h06;
      17'd12572: data = 8'h04;
      17'd12573: data = 8'h0e;
      17'd12574: data = 8'h13;
      17'd12575: data = 8'h11;
      17'd12576: data = 8'h0a;
      17'd12577: data = 8'h04;
      17'd12578: data = 8'h01;
      17'd12579: data = 8'hf5;
      17'd12580: data = 8'hf1;
      17'd12581: data = 8'hf1;
      17'd12582: data = 8'he9;
      17'd12583: data = 8'he9;
      17'd12584: data = 8'he0;
      17'd12585: data = 8'hdb;
      17'd12586: data = 8'hd6;
      17'd12587: data = 8'hd3;
      17'd12588: data = 8'hd6;
      17'd12589: data = 8'hd1;
      17'd12590: data = 8'hd5;
      17'd12591: data = 8'hda;
      17'd12592: data = 8'hdb;
      17'd12593: data = 8'hdc;
      17'd12594: data = 8'hdc;
      17'd12595: data = 8'heb;
      17'd12596: data = 8'heb;
      17'd12597: data = 8'hec;
      17'd12598: data = 8'hef;
      17'd12599: data = 8'hed;
      17'd12600: data = 8'hf5;
      17'd12601: data = 8'hf9;
      17'd12602: data = 8'hfa;
      17'd12603: data = 8'hfd;
      17'd12604: data = 8'hfd;
      17'd12605: data = 8'hfe;
      17'd12606: data = 8'h02;
      17'd12607: data = 8'hfd;
      17'd12608: data = 8'h01;
      17'd12609: data = 8'h02;
      17'd12610: data = 8'h06;
      17'd12611: data = 8'h0e;
      17'd12612: data = 8'h11;
      17'd12613: data = 8'h1a;
      17'd12614: data = 8'h1c;
      17'd12615: data = 8'h1f;
      17'd12616: data = 8'h24;
      17'd12617: data = 8'h2b;
      17'd12618: data = 8'h33;
      17'd12619: data = 8'h33;
      17'd12620: data = 8'h34;
      17'd12621: data = 8'h36;
      17'd12622: data = 8'h3a;
      17'd12623: data = 8'h3a;
      17'd12624: data = 8'h3a;
      17'd12625: data = 8'h3c;
      17'd12626: data = 8'h3c;
      17'd12627: data = 8'h39;
      17'd12628: data = 8'h33;
      17'd12629: data = 8'h2d;
      17'd12630: data = 8'h26;
      17'd12631: data = 8'h26;
      17'd12632: data = 8'h22;
      17'd12633: data = 8'h1e;
      17'd12634: data = 8'h1b;
      17'd12635: data = 8'h1a;
      17'd12636: data = 8'h1b;
      17'd12637: data = 8'h15;
      17'd12638: data = 8'h13;
      17'd12639: data = 8'h13;
      17'd12640: data = 8'h12;
      17'd12641: data = 8'h0e;
      17'd12642: data = 8'h0a;
      17'd12643: data = 8'h0d;
      17'd12644: data = 8'h0a;
      17'd12645: data = 8'h06;
      17'd12646: data = 8'h05;
      17'd12647: data = 8'h00;
      17'd12648: data = 8'hf6;
      17'd12649: data = 8'hf4;
      17'd12650: data = 8'hed;
      17'd12651: data = 8'he5;
      17'd12652: data = 8'he3;
      17'd12653: data = 8'he2;
      17'd12654: data = 8'he2;
      17'd12655: data = 8'hdb;
      17'd12656: data = 8'hd6;
      17'd12657: data = 8'hd3;
      17'd12658: data = 8'hd2;
      17'd12659: data = 8'hcd;
      17'd12660: data = 8'hca;
      17'd12661: data = 8'hcd;
      17'd12662: data = 8'hce;
      17'd12663: data = 8'hce;
      17'd12664: data = 8'hce;
      17'd12665: data = 8'hd3;
      17'd12666: data = 8'hd5;
      17'd12667: data = 8'hda;
      17'd12668: data = 8'hdc;
      17'd12669: data = 8'hdc;
      17'd12670: data = 8'hde;
      17'd12671: data = 8'he2;
      17'd12672: data = 8'he4;
      17'd12673: data = 8'he4;
      17'd12674: data = 8'he5;
      17'd12675: data = 8'heb;
      17'd12676: data = 8'heb;
      17'd12677: data = 8'he9;
      17'd12678: data = 8'he7;
      17'd12679: data = 8'he9;
      17'd12680: data = 8'he5;
      17'd12681: data = 8'he3;
      17'd12682: data = 8'he9;
      17'd12683: data = 8'heb;
      17'd12684: data = 8'hef;
      17'd12685: data = 8'hf5;
      17'd12686: data = 8'hf9;
      17'd12687: data = 8'hfc;
      17'd12688: data = 8'hfe;
      17'd12689: data = 8'h02;
      17'd12690: data = 8'h06;
      17'd12691: data = 8'h06;
      17'd12692: data = 8'h06;
      17'd12693: data = 8'h0a;
      17'd12694: data = 8'h0d;
      17'd12695: data = 8'h11;
      17'd12696: data = 8'h11;
      17'd12697: data = 8'h12;
      17'd12698: data = 8'h12;
      17'd12699: data = 8'h11;
      17'd12700: data = 8'h0e;
      17'd12701: data = 8'h09;
      17'd12702: data = 8'h05;
      17'd12703: data = 8'h01;
      17'd12704: data = 8'h01;
      17'd12705: data = 8'h00;
      17'd12706: data = 8'hfe;
      17'd12707: data = 8'h02;
      17'd12708: data = 8'hf9;
      17'd12709: data = 8'hf5;
      17'd12710: data = 8'hfc;
      17'd12711: data = 8'hfa;
      17'd12712: data = 8'hfc;
      17'd12713: data = 8'hfd;
      17'd12714: data = 8'h01;
      17'd12715: data = 8'h00;
      17'd12716: data = 8'h00;
      17'd12717: data = 8'h01;
      17'd12718: data = 8'h00;
      17'd12719: data = 8'h00;
      17'd12720: data = 8'h00;
      17'd12721: data = 8'h00;
      17'd12722: data = 8'hfe;
      17'd12723: data = 8'hfc;
      17'd12724: data = 8'hfe;
      17'd12725: data = 8'hfc;
      17'd12726: data = 8'hf9;
      17'd12727: data = 8'hfe;
      17'd12728: data = 8'hfc;
      17'd12729: data = 8'hf9;
      17'd12730: data = 8'hf9;
      17'd12731: data = 8'hf5;
      17'd12732: data = 8'hf4;
      17'd12733: data = 8'hf4;
      17'd12734: data = 8'hfe;
      17'd12735: data = 8'hfd;
      17'd12736: data = 8'h01;
      17'd12737: data = 8'h05;
      17'd12738: data = 8'h02;
      17'd12739: data = 8'h0d;
      17'd12740: data = 8'h04;
      17'd12741: data = 8'h0c;
      17'd12742: data = 8'h0e;
      17'd12743: data = 8'h06;
      17'd12744: data = 8'h12;
      17'd12745: data = 8'h11;
      17'd12746: data = 8'h0c;
      17'd12747: data = 8'h0a;
      17'd12748: data = 8'h12;
      17'd12749: data = 8'h0d;
      17'd12750: data = 8'h11;
      17'd12751: data = 8'h0c;
      17'd12752: data = 8'h0c;
      17'd12753: data = 8'h12;
      17'd12754: data = 8'h04;
      17'd12755: data = 8'h06;
      17'd12756: data = 8'h0d;
      17'd12757: data = 8'h0e;
      17'd12758: data = 8'h04;
      17'd12759: data = 8'hfe;
      17'd12760: data = 8'h02;
      17'd12761: data = 8'hfa;
      17'd12762: data = 8'hfa;
      17'd12763: data = 8'hf4;
      17'd12764: data = 8'hfc;
      17'd12765: data = 8'hfd;
      17'd12766: data = 8'hf6;
      17'd12767: data = 8'hfd;
      17'd12768: data = 8'hf5;
      17'd12769: data = 8'hfa;
      17'd12770: data = 8'hfa;
      17'd12771: data = 8'h01;
      17'd12772: data = 8'h01;
      17'd12773: data = 8'h01;
      17'd12774: data = 8'h11;
      17'd12775: data = 8'h0a;
      17'd12776: data = 8'h0a;
      17'd12777: data = 8'h0a;
      17'd12778: data = 8'h16;
      17'd12779: data = 8'h19;
      17'd12780: data = 8'h0d;
      17'd12781: data = 8'h0c;
      17'd12782: data = 8'h0c;
      17'd12783: data = 8'h06;
      17'd12784: data = 8'hfa;
      17'd12785: data = 8'h00;
      17'd12786: data = 8'h05;
      17'd12787: data = 8'h04;
      17'd12788: data = 8'h04;
      17'd12789: data = 8'h01;
      17'd12790: data = 8'h02;
      17'd12791: data = 8'hfe;
      17'd12792: data = 8'h00;
      17'd12793: data = 8'h02;
      17'd12794: data = 8'h01;
      17'd12795: data = 8'h02;
      17'd12796: data = 8'h09;
      17'd12797: data = 8'h06;
      17'd12798: data = 8'h01;
      17'd12799: data = 8'h09;
      17'd12800: data = 8'h0a;
      17'd12801: data = 8'h0d;
      17'd12802: data = 8'hfd;
      17'd12803: data = 8'hf9;
      17'd12804: data = 8'hfd;
      17'd12805: data = 8'hf1;
      17'd12806: data = 8'hed;
      17'd12807: data = 8'he9;
      17'd12808: data = 8'hed;
      17'd12809: data = 8'heb;
      17'd12810: data = 8'he0;
      17'd12811: data = 8'he0;
      17'd12812: data = 8'hda;
      17'd12813: data = 8'hd6;
      17'd12814: data = 8'hd5;
      17'd12815: data = 8'hd6;
      17'd12816: data = 8'hd8;
      17'd12817: data = 8'hd8;
      17'd12818: data = 8'hdb;
      17'd12819: data = 8'hdb;
      17'd12820: data = 8'hdb;
      17'd12821: data = 8'he3;
      17'd12822: data = 8'hec;
      17'd12823: data = 8'hf1;
      17'd12824: data = 8'hef;
      17'd12825: data = 8'hf1;
      17'd12826: data = 8'hfa;
      17'd12827: data = 8'hfc;
      17'd12828: data = 8'hfc;
      17'd12829: data = 8'h01;
      17'd12830: data = 8'h0a;
      17'd12831: data = 8'h0c;
      17'd12832: data = 8'h06;
      17'd12833: data = 8'h09;
      17'd12834: data = 8'h09;
      17'd12835: data = 8'h09;
      17'd12836: data = 8'h09;
      17'd12837: data = 8'h0e;
      17'd12838: data = 8'h15;
      17'd12839: data = 8'h1a;
      17'd12840: data = 8'h1e;
      17'd12841: data = 8'h24;
      17'd12842: data = 8'h26;
      17'd12843: data = 8'h27;
      17'd12844: data = 8'h31;
      17'd12845: data = 8'h2f;
      17'd12846: data = 8'h2f;
      17'd12847: data = 8'h31;
      17'd12848: data = 8'h35;
      17'd12849: data = 8'h3a;
      17'd12850: data = 8'h35;
      17'd12851: data = 8'h39;
      17'd12852: data = 8'h3c;
      17'd12853: data = 8'h39;
      17'd12854: data = 8'h34;
      17'd12855: data = 8'h2d;
      17'd12856: data = 8'h2c;
      17'd12857: data = 8'h27;
      17'd12858: data = 8'h22;
      17'd12859: data = 8'h1e;
      17'd12860: data = 8'h1e;
      17'd12861: data = 8'h1a;
      17'd12862: data = 8'h13;
      17'd12863: data = 8'h12;
      17'd12864: data = 8'h0c;
      17'd12865: data = 8'h0c;
      17'd12866: data = 8'h05;
      17'd12867: data = 8'h04;
      17'd12868: data = 8'h02;
      17'd12869: data = 8'h00;
      17'd12870: data = 8'h01;
      17'd12871: data = 8'hfe;
      17'd12872: data = 8'hfc;
      17'd12873: data = 8'hfc;
      17'd12874: data = 8'hfc;
      17'd12875: data = 8'hf4;
      17'd12876: data = 8'hed;
      17'd12877: data = 8'he9;
      17'd12878: data = 8'he7;
      17'd12879: data = 8'he5;
      17'd12880: data = 8'he0;
      17'd12881: data = 8'he2;
      17'd12882: data = 8'he2;
      17'd12883: data = 8'hdb;
      17'd12884: data = 8'hd8;
      17'd12885: data = 8'hd6;
      17'd12886: data = 8'hd1;
      17'd12887: data = 8'hcb;
      17'd12888: data = 8'hcb;
      17'd12889: data = 8'hce;
      17'd12890: data = 8'hce;
      17'd12891: data = 8'hce;
      17'd12892: data = 8'hd6;
      17'd12893: data = 8'hda;
      17'd12894: data = 8'hda;
      17'd12895: data = 8'hdb;
      17'd12896: data = 8'he0;
      17'd12897: data = 8'he2;
      17'd12898: data = 8'he2;
      17'd12899: data = 8'he4;
      17'd12900: data = 8'hec;
      17'd12901: data = 8'hec;
      17'd12902: data = 8'hed;
      17'd12903: data = 8'hf4;
      17'd12904: data = 8'hf6;
      17'd12905: data = 8'hf2;
      17'd12906: data = 8'hf2;
      17'd12907: data = 8'hf5;
      17'd12908: data = 8'hf1;
      17'd12909: data = 8'hf1;
      17'd12910: data = 8'hf6;
      17'd12911: data = 8'hfa;
      17'd12912: data = 8'hf5;
      17'd12913: data = 8'hf9;
      17'd12914: data = 8'h00;
      17'd12915: data = 8'h00;
      17'd12916: data = 8'hfe;
      17'd12917: data = 8'h01;
      17'd12918: data = 8'h04;
      17'd12919: data = 8'h04;
      17'd12920: data = 8'h05;
      17'd12921: data = 8'h0a;
      17'd12922: data = 8'h0d;
      17'd12923: data = 8'h0d;
      17'd12924: data = 8'h12;
      17'd12925: data = 8'h16;
      17'd12926: data = 8'h11;
      17'd12927: data = 8'h0d;
      17'd12928: data = 8'h0a;
      17'd12929: data = 8'h09;
      17'd12930: data = 8'h05;
      17'd12931: data = 8'h02;
      17'd12932: data = 8'h05;
      17'd12933: data = 8'h00;
      17'd12934: data = 8'hfc;
      17'd12935: data = 8'hfa;
      17'd12936: data = 8'hf5;
      17'd12937: data = 8'hf4;
      17'd12938: data = 8'hf5;
      17'd12939: data = 8'hf5;
      17'd12940: data = 8'hf5;
      17'd12941: data = 8'hf5;
      17'd12942: data = 8'hf6;
      17'd12943: data = 8'hfa;
      17'd12944: data = 8'hf9;
      17'd12945: data = 8'hfd;
      17'd12946: data = 8'h02;
      17'd12947: data = 8'h04;
      17'd12948: data = 8'h01;
      17'd12949: data = 8'h01;
      17'd12950: data = 8'h01;
      17'd12951: data = 8'h01;
      17'd12952: data = 8'h00;
      17'd12953: data = 8'h00;
      17'd12954: data = 8'h01;
      17'd12955: data = 8'h01;
      17'd12956: data = 8'hfa;
      17'd12957: data = 8'hfe;
      17'd12958: data = 8'hfd;
      17'd12959: data = 8'hf2;
      17'd12960: data = 8'hfe;
      17'd12961: data = 8'hfa;
      17'd12962: data = 8'hfa;
      17'd12963: data = 8'hfd;
      17'd12964: data = 8'h00;
      17'd12965: data = 8'h0a;
      17'd12966: data = 8'h04;
      17'd12967: data = 8'h0c;
      17'd12968: data = 8'h13;
      17'd12969: data = 8'h09;
      17'd12970: data = 8'h0e;
      17'd12971: data = 8'h15;
      17'd12972: data = 8'h0d;
      17'd12973: data = 8'h13;
      17'd12974: data = 8'h12;
      17'd12975: data = 8'h16;
      17'd12976: data = 8'h1b;
      17'd12977: data = 8'h0e;
      17'd12978: data = 8'h19;
      17'd12979: data = 8'h12;
      17'd12980: data = 8'h09;
      17'd12981: data = 8'h0e;
      17'd12982: data = 8'h0d;
      17'd12983: data = 8'h0c;
      17'd12984: data = 8'hfd;
      17'd12985: data = 8'hf4;
      17'd12986: data = 8'hf9;
      17'd12987: data = 8'hf6;
      17'd12988: data = 8'hef;
      17'd12989: data = 8'hf2;
      17'd12990: data = 8'h00;
      17'd12991: data = 8'hf6;
      17'd12992: data = 8'hf4;
      17'd12993: data = 8'hfc;
      17'd12994: data = 8'hfa;
      17'd12995: data = 8'hfa;
      17'd12996: data = 8'hfe;
      17'd12997: data = 8'h09;
      17'd12998: data = 8'h0c;
      17'd12999: data = 8'h02;
      17'd13000: data = 8'h0d;
      17'd13001: data = 8'h11;
      17'd13002: data = 8'h04;
      17'd13003: data = 8'h12;
      17'd13004: data = 8'h1b;
      17'd13005: data = 8'h13;
      17'd13006: data = 8'h05;
      17'd13007: data = 8'h04;
      17'd13008: data = 8'h0c;
      17'd13009: data = 8'h00;
      17'd13010: data = 8'hfa;
      17'd13011: data = 8'h0a;
      17'd13012: data = 8'h0a;
      17'd13013: data = 8'hfa;
      17'd13014: data = 8'hf6;
      17'd13015: data = 8'h01;
      17'd13016: data = 8'h00;
      17'd13017: data = 8'hfe;
      17'd13018: data = 8'h06;
      17'd13019: data = 8'h16;
      17'd13020: data = 8'h11;
      17'd13021: data = 8'h0e;
      17'd13022: data = 8'h12;
      17'd13023: data = 8'h0a;
      17'd13024: data = 8'h04;
      17'd13025: data = 8'h0c;
      17'd13026: data = 8'h13;
      17'd13027: data = 8'h0d;
      17'd13028: data = 8'h00;
      17'd13029: data = 8'h00;
      17'd13030: data = 8'hfc;
      17'd13031: data = 8'heb;
      17'd13032: data = 8'hec;
      17'd13033: data = 8'hf5;
      17'd13034: data = 8'heb;
      17'd13035: data = 8'hdc;
      17'd13036: data = 8'hd5;
      17'd13037: data = 8'hda;
      17'd13038: data = 8'hd2;
      17'd13039: data = 8'hca;
      17'd13040: data = 8'hd8;
      17'd13041: data = 8'hdc;
      17'd13042: data = 8'hd8;
      17'd13043: data = 8'hd3;
      17'd13044: data = 8'hd8;
      17'd13045: data = 8'hda;
      17'd13046: data = 8'hda;
      17'd13047: data = 8'he5;
      17'd13048: data = 8'hf1;
      17'd13049: data = 8'hf2;
      17'd13050: data = 8'hef;
      17'd13051: data = 8'hf4;
      17'd13052: data = 8'hf5;
      17'd13053: data = 8'hf4;
      17'd13054: data = 8'hfc;
      17'd13055: data = 8'h00;
      17'd13056: data = 8'hfd;
      17'd13057: data = 8'hf6;
      17'd13058: data = 8'hf5;
      17'd13059: data = 8'hfc;
      17'd13060: data = 8'hfc;
      17'd13061: data = 8'hfd;
      17'd13062: data = 8'h0d;
      17'd13063: data = 8'h15;
      17'd13064: data = 8'h16;
      17'd13065: data = 8'h16;
      17'd13066: data = 8'h1b;
      17'd13067: data = 8'h22;
      17'd13068: data = 8'h24;
      17'd13069: data = 8'h2d;
      17'd13070: data = 8'h3d;
      17'd13071: data = 8'h3c;
      17'd13072: data = 8'h3c;
      17'd13073: data = 8'h3d;
      17'd13074: data = 8'h3a;
      17'd13075: data = 8'h3c;
      17'd13076: data = 8'h3c;
      17'd13077: data = 8'h40;
      17'd13078: data = 8'h3c;
      17'd13079: data = 8'h34;
      17'd13080: data = 8'h33;
      17'd13081: data = 8'h2f;
      17'd13082: data = 8'h29;
      17'd13083: data = 8'h27;
      17'd13084: data = 8'h2b;
      17'd13085: data = 8'h23;
      17'd13086: data = 8'h1c;
      17'd13087: data = 8'h19;
      17'd13088: data = 8'h11;
      17'd13089: data = 8'h0c;
      17'd13090: data = 8'h09;
      17'd13091: data = 8'h0e;
      17'd13092: data = 8'h12;
      17'd13093: data = 8'h0c;
      17'd13094: data = 8'h0d;
      17'd13095: data = 8'h0a;
      17'd13096: data = 8'h05;
      17'd13097: data = 8'h04;
      17'd13098: data = 8'h01;
      17'd13099: data = 8'h02;
      17'd13100: data = 8'hfa;
      17'd13101: data = 8'hed;
      17'd13102: data = 8'hec;
      17'd13103: data = 8'he2;
      17'd13104: data = 8'hda;
      17'd13105: data = 8'hda;
      17'd13106: data = 8'hd8;
      17'd13107: data = 8'hd5;
      17'd13108: data = 8'hcd;
      17'd13109: data = 8'hce;
      17'd13110: data = 8'hca;
      17'd13111: data = 8'hc4;
      17'd13112: data = 8'hc9;
      17'd13113: data = 8'hcb;
      17'd13114: data = 8'hd1;
      17'd13115: data = 8'hd1;
      17'd13116: data = 8'hd1;
      17'd13117: data = 8'hd2;
      17'd13118: data = 8'hd2;
      17'd13119: data = 8'hd6;
      17'd13120: data = 8'hdc;
      17'd13121: data = 8'he2;
      17'd13122: data = 8'hde;
      17'd13123: data = 8'he2;
      17'd13124: data = 8'he5;
      17'd13125: data = 8'he3;
      17'd13126: data = 8'he5;
      17'd13127: data = 8'heb;
      17'd13128: data = 8'hec;
      17'd13129: data = 8'hed;
      17'd13130: data = 8'hed;
      17'd13131: data = 8'hed;
      17'd13132: data = 8'hed;
      17'd13133: data = 8'he9;
      17'd13134: data = 8'hf4;
      17'd13135: data = 8'hfc;
      17'd13136: data = 8'hfa;
      17'd13137: data = 8'hfd;
      17'd13138: data = 8'hfe;
      17'd13139: data = 8'h02;
      17'd13140: data = 8'h02;
      17'd13141: data = 8'h06;
      17'd13142: data = 8'h0e;
      17'd13143: data = 8'h11;
      17'd13144: data = 8'h13;
      17'd13145: data = 8'h13;
      17'd13146: data = 8'h15;
      17'd13147: data = 8'h13;
      17'd13148: data = 8'h12;
      17'd13149: data = 8'h13;
      17'd13150: data = 8'h13;
      17'd13151: data = 8'h0e;
      17'd13152: data = 8'h0d;
      17'd13153: data = 8'h09;
      17'd13154: data = 8'h01;
      17'd13155: data = 8'h00;
      17'd13156: data = 8'h01;
      17'd13157: data = 8'h01;
      17'd13158: data = 8'hfd;
      17'd13159: data = 8'hfd;
      17'd13160: data = 8'hfc;
      17'd13161: data = 8'hf9;
      17'd13162: data = 8'hf5;
      17'd13163: data = 8'hf9;
      17'd13164: data = 8'hfd;
      17'd13165: data = 8'hfc;
      17'd13166: data = 8'hfa;
      17'd13167: data = 8'hfc;
      17'd13168: data = 8'hf9;
      17'd13169: data = 8'hf6;
      17'd13170: data = 8'hfd;
      17'd13171: data = 8'h00;
      17'd13172: data = 8'hfd;
      17'd13173: data = 8'hfd;
      17'd13174: data = 8'hfd;
      17'd13175: data = 8'hf9;
      17'd13176: data = 8'hf4;
      17'd13177: data = 8'hf5;
      17'd13178: data = 8'hf6;
      17'd13179: data = 8'hf5;
      17'd13180: data = 8'hf1;
      17'd13181: data = 8'hf2;
      17'd13182: data = 8'hf4;
      17'd13183: data = 8'hec;
      17'd13184: data = 8'hf5;
      17'd13185: data = 8'hfc;
      17'd13186: data = 8'hf9;
      17'd13187: data = 8'hfd;
      17'd13188: data = 8'h02;
      17'd13189: data = 8'h04;
      17'd13190: data = 8'h01;
      17'd13191: data = 8'h01;
      17'd13192: data = 8'h11;
      17'd13193: data = 8'h0d;
      17'd13194: data = 8'h0a;
      17'd13195: data = 8'h12;
      17'd13196: data = 8'h11;
      17'd13197: data = 8'h0a;
      17'd13198: data = 8'h0e;
      17'd13199: data = 8'h12;
      17'd13200: data = 8'h11;
      17'd13201: data = 8'h12;
      17'd13202: data = 8'h0c;
      17'd13203: data = 8'h0d;
      17'd13204: data = 8'h06;
      17'd13205: data = 8'h00;
      17'd13206: data = 8'h0a;
      17'd13207: data = 8'h06;
      17'd13208: data = 8'h05;
      17'd13209: data = 8'h16;
      17'd13210: data = 8'h12;
      17'd13211: data = 8'h01;
      17'd13212: data = 8'h04;
      17'd13213: data = 8'h02;
      17'd13214: data = 8'hfe;
      17'd13215: data = 8'hf5;
      17'd13216: data = 8'hf9;
      17'd13217: data = 8'h04;
      17'd13218: data = 8'hf6;
      17'd13219: data = 8'hf6;
      17'd13220: data = 8'h05;
      17'd13221: data = 8'h00;
      17'd13222: data = 8'hf9;
      17'd13223: data = 8'h02;
      17'd13224: data = 8'h05;
      17'd13225: data = 8'hfc;
      17'd13226: data = 8'hfd;
      17'd13227: data = 8'h06;
      17'd13228: data = 8'h09;
      17'd13229: data = 8'h04;
      17'd13230: data = 8'h0d;
      17'd13231: data = 8'h1b;
      17'd13232: data = 8'h11;
      17'd13233: data = 8'h0a;
      17'd13234: data = 8'h19;
      17'd13235: data = 8'h13;
      17'd13236: data = 8'h0a;
      17'd13237: data = 8'h06;
      17'd13238: data = 8'h0d;
      17'd13239: data = 8'h0d;
      17'd13240: data = 8'h00;
      17'd13241: data = 8'h0c;
      17'd13242: data = 8'h12;
      17'd13243: data = 8'h06;
      17'd13244: data = 8'h06;
      17'd13245: data = 8'h0c;
      17'd13246: data = 8'h0c;
      17'd13247: data = 8'h05;
      17'd13248: data = 8'h02;
      17'd13249: data = 8'h0c;
      17'd13250: data = 8'h04;
      17'd13251: data = 8'h01;
      17'd13252: data = 8'h09;
      17'd13253: data = 8'h09;
      17'd13254: data = 8'h01;
      17'd13255: data = 8'hfd;
      17'd13256: data = 8'hfd;
      17'd13257: data = 8'hf6;
      17'd13258: data = 8'hef;
      17'd13259: data = 8'heb;
      17'd13260: data = 8'hed;
      17'd13261: data = 8'he7;
      17'd13262: data = 8'he0;
      17'd13263: data = 8'he4;
      17'd13264: data = 8'hdb;
      17'd13265: data = 8'hd2;
      17'd13266: data = 8'hce;
      17'd13267: data = 8'hcb;
      17'd13268: data = 8'hd1;
      17'd13269: data = 8'hd1;
      17'd13270: data = 8'hd2;
      17'd13271: data = 8'hdc;
      17'd13272: data = 8'hd8;
      17'd13273: data = 8'hd6;
      17'd13274: data = 8'he0;
      17'd13275: data = 8'he3;
      17'd13276: data = 8'he7;
      17'd13277: data = 8'he5;
      17'd13278: data = 8'hec;
      17'd13279: data = 8'hef;
      17'd13280: data = 8'hec;
      17'd13281: data = 8'hf2;
      17'd13282: data = 8'hf5;
      17'd13283: data = 8'hf6;
      17'd13284: data = 8'h00;
      17'd13285: data = 8'h05;
      17'd13286: data = 8'h04;
      17'd13287: data = 8'h01;
      17'd13288: data = 8'h02;
      17'd13289: data = 8'h09;
      17'd13290: data = 8'h0e;
      17'd13291: data = 8'h12;
      17'd13292: data = 8'h22;
      17'd13293: data = 8'h2b;
      17'd13294: data = 8'h29;
      17'd13295: data = 8'h2f;
      17'd13296: data = 8'h31;
      17'd13297: data = 8'h33;
      17'd13298: data = 8'h36;
      17'd13299: data = 8'h3a;
      17'd13300: data = 8'h40;
      17'd13301: data = 8'h3d;
      17'd13302: data = 8'h3a;
      17'd13303: data = 8'h3e;
      17'd13304: data = 8'h3d;
      17'd13305: data = 8'h3c;
      17'd13306: data = 8'h3d;
      17'd13307: data = 8'h39;
      17'd13308: data = 8'h34;
      17'd13309: data = 8'h2c;
      17'd13310: data = 8'h26;
      17'd13311: data = 8'h24;
      17'd13312: data = 8'h1e;
      17'd13313: data = 8'h1c;
      17'd13314: data = 8'h1f;
      17'd13315: data = 8'h1f;
      17'd13316: data = 8'h19;
      17'd13317: data = 8'h12;
      17'd13318: data = 8'h11;
      17'd13319: data = 8'h0a;
      17'd13320: data = 8'h04;
      17'd13321: data = 8'h04;
      17'd13322: data = 8'h05;
      17'd13323: data = 8'h00;
      17'd13324: data = 8'hf9;
      17'd13325: data = 8'hf6;
      17'd13326: data = 8'hef;
      17'd13327: data = 8'he7;
      17'd13328: data = 8'he4;
      17'd13329: data = 8'he2;
      17'd13330: data = 8'hdb;
      17'd13331: data = 8'hd3;
      17'd13332: data = 8'hce;
      17'd13333: data = 8'hcd;
      17'd13334: data = 8'hc9;
      17'd13335: data = 8'hcb;
      17'd13336: data = 8'hd1;
      17'd13337: data = 8'hca;
      17'd13338: data = 8'hcb;
      17'd13339: data = 8'hcd;
      17'd13340: data = 8'hcd;
      17'd13341: data = 8'hcb;
      17'd13342: data = 8'hce;
      17'd13343: data = 8'hd6;
      17'd13344: data = 8'hd8;
      17'd13345: data = 8'hd5;
      17'd13346: data = 8'hd6;
      17'd13347: data = 8'hda;
      17'd13348: data = 8'hd5;
      17'd13349: data = 8'hd6;
      17'd13350: data = 8'he0;
      17'd13351: data = 8'he0;
      17'd13352: data = 8'he2;
      17'd13353: data = 8'he3;
      17'd13354: data = 8'he9;
      17'd13355: data = 8'hef;
      17'd13356: data = 8'hf1;
      17'd13357: data = 8'hf9;
      17'd13358: data = 8'hfe;
      17'd13359: data = 8'hfe;
      17'd13360: data = 8'h00;
      17'd13361: data = 8'h01;
      17'd13362: data = 8'h02;
      17'd13363: data = 8'h05;
      17'd13364: data = 8'h0e;
      17'd13365: data = 8'h16;
      17'd13366: data = 8'h12;
      17'd13367: data = 8'h13;
      17'd13368: data = 8'h16;
      17'd13369: data = 8'h15;
      17'd13370: data = 8'h12;
      17'd13371: data = 8'h15;
      17'd13372: data = 8'h19;
      17'd13373: data = 8'h15;
      17'd13374: data = 8'h11;
      17'd13375: data = 8'h11;
      17'd13376: data = 8'h13;
      17'd13377: data = 8'h0d;
      17'd13378: data = 8'h0e;
      17'd13379: data = 8'h12;
      17'd13380: data = 8'h0d;
      17'd13381: data = 8'h06;
      17'd13382: data = 8'h05;
      17'd13383: data = 8'h05;
      17'd13384: data = 8'h02;
      17'd13385: data = 8'h02;
      17'd13386: data = 8'h05;
      17'd13387: data = 8'h04;
      17'd13388: data = 8'hfd;
      17'd13389: data = 8'hf9;
      17'd13390: data = 8'hf9;
      17'd13391: data = 8'hf2;
      17'd13392: data = 8'hf1;
      17'd13393: data = 8'hf4;
      17'd13394: data = 8'hf1;
      17'd13395: data = 8'hef;
      17'd13396: data = 8'hec;
      17'd13397: data = 8'hec;
      17'd13398: data = 8'he9;
      17'd13399: data = 8'he7;
      17'd13400: data = 8'hec;
      17'd13401: data = 8'hf1;
      17'd13402: data = 8'hef;
      17'd13403: data = 8'hef;
      17'd13404: data = 8'hf2;
      17'd13405: data = 8'hf1;
      17'd13406: data = 8'hf1;
      17'd13407: data = 8'hf5;
      17'd13408: data = 8'hf9;
      17'd13409: data = 8'hfc;
      17'd13410: data = 8'hf9;
      17'd13411: data = 8'hfa;
      17'd13412: data = 8'hfd;
      17'd13413: data = 8'hf5;
      17'd13414: data = 8'h02;
      17'd13415: data = 8'h05;
      17'd13416: data = 8'hfc;
      17'd13417: data = 8'h0c;
      17'd13418: data = 8'h05;
      17'd13419: data = 8'h04;
      17'd13420: data = 8'h0e;
      17'd13421: data = 8'h04;
      17'd13422: data = 8'h11;
      17'd13423: data = 8'h19;
      17'd13424: data = 8'h0c;
      17'd13425: data = 8'h15;
      17'd13426: data = 8'h12;
      17'd13427: data = 8'h09;
      17'd13428: data = 8'h19;
      17'd13429: data = 8'h16;
      17'd13430: data = 8'h11;
      17'd13431: data = 8'h1f;
      17'd13432: data = 8'h19;
      17'd13433: data = 8'h12;
      17'd13434: data = 8'h15;
      17'd13435: data = 8'h0e;
      17'd13436: data = 8'h0d;
      17'd13437: data = 8'h06;
      17'd13438: data = 8'hfe;
      17'd13439: data = 8'h01;
      17'd13440: data = 8'hfa;
      17'd13441: data = 8'heb;
      17'd13442: data = 8'hef;
      17'd13443: data = 8'he9;
      17'd13444: data = 8'he5;
      17'd13445: data = 8'hfe;
      17'd13446: data = 8'h00;
      17'd13447: data = 8'h04;
      17'd13448: data = 8'h0e;
      17'd13449: data = 8'h16;
      17'd13450: data = 8'h1f;
      17'd13451: data = 8'h16;
      17'd13452: data = 8'h11;
      17'd13453: data = 8'h1b;
      17'd13454: data = 8'h12;
      17'd13455: data = 8'h0d;
      17'd13456: data = 8'h19;
      17'd13457: data = 8'h13;
      17'd13458: data = 8'h0a;
      17'd13459: data = 8'h09;
      17'd13460: data = 8'h01;
      17'd13461: data = 8'h02;
      17'd13462: data = 8'hfa;
      17'd13463: data = 8'hf6;
      17'd13464: data = 8'h00;
      17'd13465: data = 8'hf2;
      17'd13466: data = 8'hfc;
      17'd13467: data = 8'h0d;
      17'd13468: data = 8'h0d;
      17'd13469: data = 8'h15;
      17'd13470: data = 8'h1f;
      17'd13471: data = 8'h26;
      17'd13472: data = 8'h22;
      17'd13473: data = 8'h11;
      17'd13474: data = 8'h12;
      17'd13475: data = 8'h12;
      17'd13476: data = 8'h06;
      17'd13477: data = 8'h09;
      17'd13478: data = 8'h09;
      17'd13479: data = 8'hfe;
      17'd13480: data = 8'hf2;
      17'd13481: data = 8'he4;
      17'd13482: data = 8'hdc;
      17'd13483: data = 8'hd6;
      17'd13484: data = 8'hd1;
      17'd13485: data = 8'hd6;
      17'd13486: data = 8'hd3;
      17'd13487: data = 8'hcd;
      17'd13488: data = 8'hd3;
      17'd13489: data = 8'hdb;
      17'd13490: data = 8'hda;
      17'd13491: data = 8'he2;
      17'd13492: data = 8'hec;
      17'd13493: data = 8'hec;
      17'd13494: data = 8'he9;
      17'd13495: data = 8'hdb;
      17'd13496: data = 8'hde;
      17'd13497: data = 8'hdc;
      17'd13498: data = 8'hd6;
      17'd13499: data = 8'he2;
      17'd13500: data = 8'he2;
      17'd13501: data = 8'hdb;
      17'd13502: data = 8'hd5;
      17'd13503: data = 8'hcd;
      17'd13504: data = 8'hce;
      17'd13505: data = 8'hd5;
      17'd13506: data = 8'he0;
      17'd13507: data = 8'hef;
      17'd13508: data = 8'hf6;
      17'd13509: data = 8'hfc;
      17'd13510: data = 8'h09;
      17'd13511: data = 8'h11;
      17'd13512: data = 8'h16;
      17'd13513: data = 8'h23;
      17'd13514: data = 8'h2b;
      17'd13515: data = 8'h31;
      17'd13516: data = 8'h29;
      17'd13517: data = 8'h26;
      17'd13518: data = 8'h2b;
      17'd13519: data = 8'h27;
      17'd13520: data = 8'h2c;
      17'd13521: data = 8'h35;
      17'd13522: data = 8'h33;
      17'd13523: data = 8'h2d;
      17'd13524: data = 8'h2b;
      17'd13525: data = 8'h24;
      17'd13526: data = 8'h24;
      17'd13527: data = 8'h2b;
      17'd13528: data = 8'h34;
      17'd13529: data = 8'h3e;
      17'd13530: data = 8'h3c;
      17'd13531: data = 8'h40;
      17'd13532: data = 8'h43;
      17'd13533: data = 8'h3d;
      17'd13534: data = 8'h3e;
      17'd13535: data = 8'h3c;
      17'd13536: data = 8'h3a;
      17'd13537: data = 8'h33;
      17'd13538: data = 8'h24;
      17'd13539: data = 8'h1c;
      17'd13540: data = 8'h13;
      17'd13541: data = 8'h0d;
      17'd13542: data = 8'h0c;
      17'd13543: data = 8'h0a;
      17'd13544: data = 8'h00;
      17'd13545: data = 8'hf9;
      17'd13546: data = 8'hed;
      17'd13547: data = 8'he3;
      17'd13548: data = 8'he3;
      17'd13549: data = 8'he4;
      17'd13550: data = 8'hed;
      17'd13551: data = 8'hf4;
      17'd13552: data = 8'hef;
      17'd13553: data = 8'hef;
      17'd13554: data = 8'he9;
      17'd13555: data = 8'he2;
      17'd13556: data = 8'he2;
      17'd13557: data = 8'he2;
      17'd13558: data = 8'he0;
      17'd13559: data = 8'hd8;
      17'd13560: data = 8'hd1;
      17'd13561: data = 8'hcb;
      17'd13562: data = 8'hc9;
      17'd13563: data = 8'hc5;
      17'd13564: data = 8'hc9;
      17'd13565: data = 8'hc6;
      17'd13566: data = 8'hc4;
      17'd13567: data = 8'hc2;
      17'd13568: data = 8'hc1;
      17'd13569: data = 8'hc6;
      17'd13570: data = 8'hcd;
      17'd13571: data = 8'hdc;
      17'd13572: data = 8'he9;
      17'd13573: data = 8'hec;
      17'd13574: data = 8'hf1;
      17'd13575: data = 8'hf4;
      17'd13576: data = 8'hf1;
      17'd13577: data = 8'hed;
      17'd13578: data = 8'hef;
      17'd13579: data = 8'hf4;
      17'd13580: data = 8'hf9;
      17'd13581: data = 8'hf9;
      17'd13582: data = 8'hfa;
      17'd13583: data = 8'hfc;
      17'd13584: data = 8'hfa;
      17'd13585: data = 8'h01;
      17'd13586: data = 8'h09;
      17'd13587: data = 8'h06;
      17'd13588: data = 8'h06;
      17'd13589: data = 8'h09;
      17'd13590: data = 8'h0c;
      17'd13591: data = 8'h11;
      17'd13592: data = 8'h1a;
      17'd13593: data = 8'h22;
      17'd13594: data = 8'h24;
      17'd13595: data = 8'h23;
      17'd13596: data = 8'h22;
      17'd13597: data = 8'h1f;
      17'd13598: data = 8'h15;
      17'd13599: data = 8'h12;
      17'd13600: data = 8'h11;
      17'd13601: data = 8'h0d;
      17'd13602: data = 8'h0a;
      17'd13603: data = 8'h05;
      17'd13604: data = 8'h02;
      17'd13605: data = 8'h00;
      17'd13606: data = 8'h00;
      17'd13607: data = 8'hfe;
      17'd13608: data = 8'hfc;
      17'd13609: data = 8'hf9;
      17'd13610: data = 8'hf6;
      17'd13611: data = 8'hf5;
      17'd13612: data = 8'hf4;
      17'd13613: data = 8'hf6;
      17'd13614: data = 8'hfd;
      17'd13615: data = 8'hfe;
      17'd13616: data = 8'hfc;
      17'd13617: data = 8'hf4;
      17'd13618: data = 8'hef;
      17'd13619: data = 8'he7;
      17'd13620: data = 8'he0;
      17'd13621: data = 8'he0;
      17'd13622: data = 8'he0;
      17'd13623: data = 8'he3;
      17'd13624: data = 8'he5;
      17'd13625: data = 8'he4;
      17'd13626: data = 8'he4;
      17'd13627: data = 8'he5;
      17'd13628: data = 8'hec;
      17'd13629: data = 8'hef;
      17'd13630: data = 8'hf2;
      17'd13631: data = 8'hf6;
      17'd13632: data = 8'hf5;
      17'd13633: data = 8'hf9;
      17'd13634: data = 8'hfa;
      17'd13635: data = 8'hfe;
      17'd13636: data = 8'h06;
      17'd13637: data = 8'h05;
      17'd13638: data = 8'h04;
      17'd13639: data = 8'h04;
      17'd13640: data = 8'hfa;
      17'd13641: data = 8'hfd;
      17'd13642: data = 8'h02;
      17'd13643: data = 8'hfe;
      17'd13644: data = 8'h0a;
      17'd13645: data = 8'h16;
      17'd13646: data = 8'h0c;
      17'd13647: data = 8'h1a;
      17'd13648: data = 8'h1c;
      17'd13649: data = 8'h0c;
      17'd13650: data = 8'h22;
      17'd13651: data = 8'h1a;
      17'd13652: data = 8'h15;
      17'd13653: data = 8'h24;
      17'd13654: data = 8'h11;
      17'd13655: data = 8'h12;
      17'd13656: data = 8'h1c;
      17'd13657: data = 8'h0c;
      17'd13658: data = 8'h12;
      17'd13659: data = 8'h1b;
      17'd13660: data = 8'h09;
      17'd13661: data = 8'h02;
      17'd13662: data = 8'h01;
      17'd13663: data = 8'hf5;
      17'd13664: data = 8'hfd;
      17'd13665: data = 8'hf6;
      17'd13666: data = 8'h02;
      17'd13667: data = 8'h0a;
      17'd13668: data = 8'hed;
      17'd13669: data = 8'hf1;
      17'd13670: data = 8'h02;
      17'd13671: data = 8'hf2;
      17'd13672: data = 8'hf6;
      17'd13673: data = 8'h1a;
      17'd13674: data = 8'h1b;
      17'd13675: data = 8'h1f;
      17'd13676: data = 8'h16;
      17'd13677: data = 8'h0d;
      17'd13678: data = 8'h12;
      17'd13679: data = 8'hf2;
      17'd13680: data = 8'h01;
      17'd13681: data = 8'h12;
      17'd13682: data = 8'hfc;
      17'd13683: data = 8'hfa;
      17'd13684: data = 8'hfa;
      17'd13685: data = 8'hf9;
      17'd13686: data = 8'hf5;
      17'd13687: data = 8'h02;
      17'd13688: data = 8'h1b;
      17'd13689: data = 8'h1c;
      17'd13690: data = 8'h0d;
      17'd13691: data = 8'h19;
      17'd13692: data = 8'h1f;
      17'd13693: data = 8'h04;
      17'd13694: data = 8'h13;
      17'd13695: data = 8'h27;
      17'd13696: data = 8'h2c;
      17'd13697: data = 8'h22;
      17'd13698: data = 8'h0a;
      17'd13699: data = 8'h01;
      17'd13700: data = 8'heb;
      17'd13701: data = 8'he2;
      17'd13702: data = 8'hf1;
      17'd13703: data = 8'hf4;
      17'd13704: data = 8'hf2;
      17'd13705: data = 8'hf5;
      17'd13706: data = 8'hed;
      17'd13707: data = 8'he5;
      17'd13708: data = 8'he7;
      17'd13709: data = 8'hf1;
      17'd13710: data = 8'h04;
      17'd13711: data = 8'hfc;
      17'd13712: data = 8'hf1;
      17'd13713: data = 8'hec;
      17'd13714: data = 8'hd1;
      17'd13715: data = 8'hc9;
      17'd13716: data = 8'hd2;
      17'd13717: data = 8'hda;
      17'd13718: data = 8'hdb;
      17'd13719: data = 8'hd6;
      17'd13720: data = 8'hc6;
      17'd13721: data = 8'hbb;
      17'd13722: data = 8'hb5;
      17'd13723: data = 8'hc1;
      17'd13724: data = 8'hda;
      17'd13725: data = 8'he0;
      17'd13726: data = 8'hf4;
      17'd13727: data = 8'hfa;
      17'd13728: data = 8'heb;
      17'd13729: data = 8'hf2;
      17'd13730: data = 8'hf4;
      17'd13731: data = 8'hfe;
      17'd13732: data = 8'h0c;
      17'd13733: data = 8'h06;
      17'd13734: data = 8'h05;
      17'd13735: data = 8'hfc;
      17'd13736: data = 8'hf1;
      17'd13737: data = 8'hfa;
      17'd13738: data = 8'h09;
      17'd13739: data = 8'h13;
      17'd13740: data = 8'h29;
      17'd13741: data = 8'h29;
      17'd13742: data = 8'h1e;
      17'd13743: data = 8'h1e;
      17'd13744: data = 8'h23;
      17'd13745: data = 8'h35;
      17'd13746: data = 8'h43;
      17'd13747: data = 8'h52;
      17'd13748: data = 8'h5c;
      17'd13749: data = 8'h4e;
      17'd13750: data = 8'h3e;
      17'd13751: data = 8'h3c;
      17'd13752: data = 8'h34;
      17'd13753: data = 8'h34;
      17'd13754: data = 8'h39;
      17'd13755: data = 8'h31;
      17'd13756: data = 8'h2b;
      17'd13757: data = 8'h1f;
      17'd13758: data = 8'h1a;
      17'd13759: data = 8'h26;
      17'd13760: data = 8'h27;
      17'd13761: data = 8'h34;
      17'd13762: data = 8'h39;
      17'd13763: data = 8'h2c;
      17'd13764: data = 8'h22;
      17'd13765: data = 8'h19;
      17'd13766: data = 8'h13;
      17'd13767: data = 8'h11;
      17'd13768: data = 8'h0d;
      17'd13769: data = 8'h0e;
      17'd13770: data = 8'h0c;
      17'd13771: data = 8'hf4;
      17'd13772: data = 8'he2;
      17'd13773: data = 8'hdc;
      17'd13774: data = 8'hd2;
      17'd13775: data = 8'hd6;
      17'd13776: data = 8'hdc;
      17'd13777: data = 8'hd6;
      17'd13778: data = 8'hda;
      17'd13779: data = 8'hd5;
      17'd13780: data = 8'hd6;
      17'd13781: data = 8'hdc;
      17'd13782: data = 8'hde;
      17'd13783: data = 8'he9;
      17'd13784: data = 8'he7;
      17'd13785: data = 8'hda;
      17'd13786: data = 8'hd1;
      17'd13787: data = 8'hc6;
      17'd13788: data = 8'hc5;
      17'd13789: data = 8'hc9;
      17'd13790: data = 8'hca;
      17'd13791: data = 8'hd1;
      17'd13792: data = 8'hcd;
      17'd13793: data = 8'hc5;
      17'd13794: data = 8'hc6;
      17'd13795: data = 8'hcd;
      17'd13796: data = 8'hd5;
      17'd13797: data = 8'he3;
      17'd13798: data = 8'hec;
      17'd13799: data = 8'hf2;
      17'd13800: data = 8'hf6;
      17'd13801: data = 8'hf9;
      17'd13802: data = 8'hf6;
      17'd13803: data = 8'hfd;
      17'd13804: data = 8'h02;
      17'd13805: data = 8'h0a;
      17'd13806: data = 8'h04;
      17'd13807: data = 8'hfc;
      17'd13808: data = 8'hfa;
      17'd13809: data = 8'hf6;
      17'd13810: data = 8'hfe;
      17'd13811: data = 8'h0a;
      17'd13812: data = 8'h11;
      17'd13813: data = 8'h19;
      17'd13814: data = 8'h1e;
      17'd13815: data = 8'h1b;
      17'd13816: data = 8'h1b;
      17'd13817: data = 8'h1b;
      17'd13818: data = 8'h1f;
      17'd13819: data = 8'h29;
      17'd13820: data = 8'h26;
      17'd13821: data = 8'h1e;
      17'd13822: data = 8'h1c;
      17'd13823: data = 8'h12;
      17'd13824: data = 8'h0a;
      17'd13825: data = 8'h09;
      17'd13826: data = 8'h0a;
      17'd13827: data = 8'h09;
      17'd13828: data = 8'h01;
      17'd13829: data = 8'hfa;
      17'd13830: data = 8'hf9;
      17'd13831: data = 8'hf6;
      17'd13832: data = 8'hfa;
      17'd13833: data = 8'h02;
      17'd13834: data = 8'h02;
      17'd13835: data = 8'h01;
      17'd13836: data = 8'hfc;
      17'd13837: data = 8'hf1;
      17'd13838: data = 8'heb;
      17'd13839: data = 8'he5;
      17'd13840: data = 8'heb;
      17'd13841: data = 8'hec;
      17'd13842: data = 8'he5;
      17'd13843: data = 8'he0;
      17'd13844: data = 8'hde;
      17'd13845: data = 8'hdb;
      17'd13846: data = 8'hda;
      17'd13847: data = 8'hdc;
      17'd13848: data = 8'he5;
      17'd13849: data = 8'he7;
      17'd13850: data = 8'he3;
      17'd13851: data = 8'he3;
      17'd13852: data = 8'he7;
      17'd13853: data = 8'he9;
      17'd13854: data = 8'hf1;
      17'd13855: data = 8'hfc;
      17'd13856: data = 8'hfc;
      17'd13857: data = 8'hfd;
      17'd13858: data = 8'hf9;
      17'd13859: data = 8'hf1;
      17'd13860: data = 8'hf2;
      17'd13861: data = 8'hf9;
      17'd13862: data = 8'h04;
      17'd13863: data = 8'h0c;
      17'd13864: data = 8'h05;
      17'd13865: data = 8'h0c;
      17'd13866: data = 8'h0d;
      17'd13867: data = 8'h0c;
      17'd13868: data = 8'h13;
      17'd13869: data = 8'h15;
      17'd13870: data = 8'h16;
      17'd13871: data = 8'h1c;
      17'd13872: data = 8'h15;
      17'd13873: data = 8'h0e;
      17'd13874: data = 8'h13;
      17'd13875: data = 8'h16;
      17'd13876: data = 8'h1b;
      17'd13877: data = 8'h16;
      17'd13878: data = 8'h16;
      17'd13879: data = 8'h1c;
      17'd13880: data = 8'h11;
      17'd13881: data = 8'h11;
      17'd13882: data = 8'h16;
      17'd13883: data = 8'h1b;
      17'd13884: data = 8'h1e;
      17'd13885: data = 8'h1c;
      17'd13886: data = 8'h1a;
      17'd13887: data = 8'h0c;
      17'd13888: data = 8'h00;
      17'd13889: data = 8'hf6;
      17'd13890: data = 8'hf2;
      17'd13891: data = 8'hec;
      17'd13892: data = 8'hec;
      17'd13893: data = 8'hfa;
      17'd13894: data = 8'hef;
      17'd13895: data = 8'hef;
      17'd13896: data = 8'hf6;
      17'd13897: data = 8'hfe;
      17'd13898: data = 8'hf9;
      17'd13899: data = 8'hf9;
      17'd13900: data = 8'h05;
      17'd13901: data = 8'h06;
      17'd13902: data = 8'h02;
      17'd13903: data = 8'h04;
      17'd13904: data = 8'h0e;
      17'd13905: data = 8'h0a;
      17'd13906: data = 8'h02;
      17'd13907: data = 8'h02;
      17'd13908: data = 8'hfa;
      17'd13909: data = 8'hf6;
      17'd13910: data = 8'hf4;
      17'd13911: data = 8'hf9;
      17'd13912: data = 8'hfc;
      17'd13913: data = 8'hfd;
      17'd13914: data = 8'h0e;
      17'd13915: data = 8'h1a;
      17'd13916: data = 8'h1b;
      17'd13917: data = 8'h22;
      17'd13918: data = 8'h29;
      17'd13919: data = 8'h1b;
      17'd13920: data = 8'h13;
      17'd13921: data = 8'h12;
      17'd13922: data = 8'h0e;
      17'd13923: data = 8'h09;
      17'd13924: data = 8'h02;
      17'd13925: data = 8'h09;
      17'd13926: data = 8'h01;
      17'd13927: data = 8'hfe;
      17'd13928: data = 8'h00;
      17'd13929: data = 8'hfa;
      17'd13930: data = 8'hfc;
      17'd13931: data = 8'hfd;
      17'd13932: data = 8'hfe;
      17'd13933: data = 8'hfa;
      17'd13934: data = 8'hf9;
      17'd13935: data = 8'hf9;
      17'd13936: data = 8'hf6;
      17'd13937: data = 8'hec;
      17'd13938: data = 8'he5;
      17'd13939: data = 8'he3;
      17'd13940: data = 8'hd5;
      17'd13941: data = 8'hca;
      17'd13942: data = 8'hc5;
      17'd13943: data = 8'hc4;
      17'd13944: data = 8'hc9;
      17'd13945: data = 8'hcb;
      17'd13946: data = 8'hd6;
      17'd13947: data = 8'hdc;
      17'd13948: data = 8'hdb;
      17'd13949: data = 8'he0;
      17'd13950: data = 8'hde;
      17'd13951: data = 8'hdc;
      17'd13952: data = 8'he0;
      17'd13953: data = 8'he3;
      17'd13954: data = 8'he0;
      17'd13955: data = 8'he0;
      17'd13956: data = 8'he3;
      17'd13957: data = 8'he5;
      17'd13958: data = 8'hec;
      17'd13959: data = 8'hef;
      17'd13960: data = 8'hf9;
      17'd13961: data = 8'hfe;
      17'd13962: data = 8'h01;
      17'd13963: data = 8'h09;
      17'd13964: data = 8'h0e;
      17'd13965: data = 8'h16;
      17'd13966: data = 8'h1f;
      17'd13967: data = 8'h29;
      17'd13968: data = 8'h2d;
      17'd13969: data = 8'h2f;
      17'd13970: data = 8'h2d;
      17'd13971: data = 8'h2c;
      17'd13972: data = 8'h29;
      17'd13973: data = 8'h27;
      17'd13974: data = 8'h31;
      17'd13975: data = 8'h33;
      17'd13976: data = 8'h34;
      17'd13977: data = 8'h3d;
      17'd13978: data = 8'h40;
      17'd13979: data = 8'h43;
      17'd13980: data = 8'h40;
      17'd13981: data = 8'h40;
      17'd13982: data = 8'h3e;
      17'd13983: data = 8'h36;
      17'd13984: data = 8'h33;
      17'd13985: data = 8'h2c;
      17'd13986: data = 8'h26;
      17'd13987: data = 8'h22;
      17'd13988: data = 8'h24;
      17'd13989: data = 8'h23;
      17'd13990: data = 8'h1c;
      17'd13991: data = 8'h19;
      17'd13992: data = 8'h12;
      17'd13993: data = 8'h0a;
      17'd13994: data = 8'h04;
      17'd13995: data = 8'h04;
      17'd13996: data = 8'h02;
      17'd13997: data = 8'hfd;
      17'd13998: data = 8'hf9;
      17'd13999: data = 8'hf6;
      17'd14000: data = 8'hef;
      17'd14001: data = 8'he3;
      17'd14002: data = 8'hda;
      17'd14003: data = 8'hd6;
      17'd14004: data = 8'hd2;
      17'd14005: data = 8'hca;
      17'd14006: data = 8'hca;
      17'd14007: data = 8'hce;
      17'd14008: data = 8'hd2;
      17'd14009: data = 8'hd5;
      17'd14010: data = 8'hd8;
      17'd14011: data = 8'hd8;
      17'd14012: data = 8'hd6;
      17'd14013: data = 8'hd5;
      17'd14014: data = 8'hce;
      17'd14015: data = 8'hca;
      17'd14016: data = 8'hc9;
      17'd14017: data = 8'hca;
      17'd14018: data = 8'hcd;
      17'd14019: data = 8'hce;
      17'd14020: data = 8'hd3;
      17'd14021: data = 8'hd8;
      17'd14022: data = 8'hdc;
      17'd14023: data = 8'hda;
      17'd14024: data = 8'hdb;
      17'd14025: data = 8'heb;
      17'd14026: data = 8'hec;
      17'd14027: data = 8'heb;
      17'd14028: data = 8'hf5;
      17'd14029: data = 8'h02;
      17'd14030: data = 8'h04;
      17'd14031: data = 8'h01;
      17'd14032: data = 8'h02;
      17'd14033: data = 8'h02;
      17'd14034: data = 8'h02;
      17'd14035: data = 8'h04;
      17'd14036: data = 8'h04;
      17'd14037: data = 8'h05;
      17'd14038: data = 8'h0e;
      17'd14039: data = 8'h1a;
      17'd14040: data = 8'h1e;
      17'd14041: data = 8'h22;
      17'd14042: data = 8'h23;
      17'd14043: data = 8'h24;
      17'd14044: data = 8'h1f;
      17'd14045: data = 8'h1a;
      17'd14046: data = 8'h1c;
      17'd14047: data = 8'h1a;
      17'd14048: data = 8'h12;
      17'd14049: data = 8'h0d;
      17'd14050: data = 8'h15;
      17'd14051: data = 8'h12;
      17'd14052: data = 8'h0c;
      17'd14053: data = 8'h0a;
      17'd14054: data = 8'h09;
      17'd14055: data = 8'h09;
      17'd14056: data = 8'h05;
      17'd14057: data = 8'h01;
      17'd14058: data = 8'hfe;
      17'd14059: data = 8'hfe;
      17'd14060: data = 8'h02;
      17'd14061: data = 8'hfd;
      17'd14062: data = 8'hf2;
      17'd14063: data = 8'hec;
      17'd14064: data = 8'he5;
      17'd14065: data = 8'he4;
      17'd14066: data = 8'he0;
      17'd14067: data = 8'hdb;
      17'd14068: data = 8'he2;
      17'd14069: data = 8'he7;
      17'd14070: data = 8'he9;
      17'd14071: data = 8'hec;
      17'd14072: data = 8'hf1;
      17'd14073: data = 8'hec;
      17'd14074: data = 8'he9;
      17'd14075: data = 8'he4;
      17'd14076: data = 8'he2;
      17'd14077: data = 8'he2;
      17'd14078: data = 8'he0;
      17'd14079: data = 8'he0;
      17'd14080: data = 8'he4;
      17'd14081: data = 8'hef;
      17'd14082: data = 8'hf5;
      17'd14083: data = 8'hf2;
      17'd14084: data = 8'hfd;
      17'd14085: data = 8'h01;
      17'd14086: data = 8'h02;
      17'd14087: data = 8'h01;
      17'd14088: data = 8'hfd;
      17'd14089: data = 8'h05;
      17'd14090: data = 8'h0d;
      17'd14091: data = 8'h09;
      17'd14092: data = 8'h12;
      17'd14093: data = 8'h11;
      17'd14094: data = 8'hf6;
      17'd14095: data = 8'h09;
      17'd14096: data = 8'h1a;
      17'd14097: data = 8'h1b;
      17'd14098: data = 8'h15;
      17'd14099: data = 8'h1e;
      17'd14100: data = 8'h1a;
      17'd14101: data = 8'h11;
      17'd14102: data = 8'h23;
      17'd14103: data = 8'h23;
      17'd14104: data = 8'h1b;
      17'd14105: data = 8'h1a;
      17'd14106: data = 8'h12;
      17'd14107: data = 8'h09;
      17'd14108: data = 8'h0d;
      17'd14109: data = 8'h12;
      17'd14110: data = 8'h06;
      17'd14111: data = 8'h12;
      17'd14112: data = 8'h1f;
      17'd14113: data = 8'h13;
      17'd14114: data = 8'h16;
      17'd14115: data = 8'h11;
      17'd14116: data = 8'h06;
      17'd14117: data = 8'h00;
      17'd14118: data = 8'hf2;
      17'd14119: data = 8'hf5;
      17'd14120: data = 8'hf1;
      17'd14121: data = 8'hf4;
      17'd14122: data = 8'hfd;
      17'd14123: data = 8'hed;
      17'd14124: data = 8'hdc;
      17'd14125: data = 8'hd8;
      17'd14126: data = 8'hef;
      17'd14127: data = 8'h09;
      17'd14128: data = 8'h00;
      17'd14129: data = 8'h11;
      17'd14130: data = 8'h31;
      17'd14131: data = 8'h33;
      17'd14132: data = 8'h12;
      17'd14133: data = 8'hf6;
      17'd14134: data = 8'he5;
      17'd14135: data = 8'hd3;
      17'd14136: data = 8'hd8;
      17'd14137: data = 8'he5;
      17'd14138: data = 8'hfa;
      17'd14139: data = 8'h06;
      17'd14140: data = 8'h0e;
      17'd14141: data = 8'h1b;
      17'd14142: data = 8'h23;
      17'd14143: data = 8'h2c;
      17'd14144: data = 8'h34;
      17'd14145: data = 8'h2f;
      17'd14146: data = 8'h19;
      17'd14147: data = 8'hfd;
      17'd14148: data = 8'hf6;
      17'd14149: data = 8'hef;
      17'd14150: data = 8'hef;
      17'd14151: data = 8'h13;
      17'd14152: data = 8'h33;
      17'd14153: data = 8'h1f;
      17'd14154: data = 8'hfa;
      17'd14155: data = 8'hf6;
      17'd14156: data = 8'h00;
      17'd14157: data = 8'h02;
      17'd14158: data = 8'h12;
      17'd14159: data = 8'h22;
      17'd14160: data = 8'h22;
      17'd14161: data = 8'h19;
      17'd14162: data = 8'h01;
      17'd14163: data = 8'he0;
      17'd14164: data = 8'hca;
      17'd14165: data = 8'hd3;
      17'd14166: data = 8'he2;
      17'd14167: data = 8'he0;
      17'd14168: data = 8'hdb;
      17'd14169: data = 8'hd8;
      17'd14170: data = 8'he2;
      17'd14171: data = 8'he7;
      17'd14172: data = 8'hec;
      17'd14173: data = 8'hfa;
      17'd14174: data = 8'hfd;
      17'd14175: data = 8'hdc;
      17'd14176: data = 8'hc5;
      17'd14177: data = 8'hbd;
      17'd14178: data = 8'hb5;
      17'd14179: data = 8'hc0;
      17'd14180: data = 8'hd6;
      17'd14181: data = 8'hf1;
      17'd14182: data = 8'hf5;
      17'd14183: data = 8'hf1;
      17'd14184: data = 8'he0;
      17'd14185: data = 8'hd5;
      17'd14186: data = 8'he5;
      17'd14187: data = 8'hfa;
      17'd14188: data = 8'h00;
      17'd14189: data = 8'h00;
      17'd14190: data = 8'h01;
      17'd14191: data = 8'h06;
      17'd14192: data = 8'h06;
      17'd14193: data = 8'h02;
      17'd14194: data = 8'h05;
      17'd14195: data = 8'h12;
      17'd14196: data = 8'h1c;
      17'd14197: data = 8'h15;
      17'd14198: data = 8'h12;
      17'd14199: data = 8'h1a;
      17'd14200: data = 8'h2b;
      17'd14201: data = 8'h3d;
      17'd14202: data = 8'h45;
      17'd14203: data = 8'h47;
      17'd14204: data = 8'h40;
      17'd14205: data = 8'h33;
      17'd14206: data = 8'h26;
      17'd14207: data = 8'h1a;
      17'd14208: data = 8'h22;
      17'd14209: data = 8'h29;
      17'd14210: data = 8'h2f;
      17'd14211: data = 8'h3c;
      17'd14212: data = 8'h40;
      17'd14213: data = 8'h3d;
      17'd14214: data = 8'h33;
      17'd14215: data = 8'h29;
      17'd14216: data = 8'h29;
      17'd14217: data = 8'h27;
      17'd14218: data = 8'h24;
      17'd14219: data = 8'h13;
      17'd14220: data = 8'h0a;
      17'd14221: data = 8'h11;
      17'd14222: data = 8'h0e;
      17'd14223: data = 8'h09;
      17'd14224: data = 8'h01;
      17'd14225: data = 8'h00;
      17'd14226: data = 8'hfe;
      17'd14227: data = 8'hf4;
      17'd14228: data = 8'he5;
      17'd14229: data = 8'he3;
      17'd14230: data = 8'hed;
      17'd14231: data = 8'hf4;
      17'd14232: data = 8'hf2;
      17'd14233: data = 8'hef;
      17'd14234: data = 8'he3;
      17'd14235: data = 8'hd8;
      17'd14236: data = 8'hcd;
      17'd14237: data = 8'hc5;
      17'd14238: data = 8'hca;
      17'd14239: data = 8'hd5;
      17'd14240: data = 8'hd6;
      17'd14241: data = 8'hda;
      17'd14242: data = 8'hde;
      17'd14243: data = 8'hde;
      17'd14244: data = 8'hda;
      17'd14245: data = 8'hd6;
      17'd14246: data = 8'hd5;
      17'd14247: data = 8'hd5;
      17'd14248: data = 8'hd1;
      17'd14249: data = 8'hca;
      17'd14250: data = 8'hcb;
      17'd14251: data = 8'hd8;
      17'd14252: data = 8'he7;
      17'd14253: data = 8'hef;
      17'd14254: data = 8'heb;
      17'd14255: data = 8'he9;
      17'd14256: data = 8'hed;
      17'd14257: data = 8'hec;
      17'd14258: data = 8'heb;
      17'd14259: data = 8'hf4;
      17'd14260: data = 8'hfe;
      17'd14261: data = 8'h05;
      17'd14262: data = 8'h0d;
      17'd14263: data = 8'h0d;
      17'd14264: data = 8'h0a;
      17'd14265: data = 8'h06;
      17'd14266: data = 8'h04;
      17'd14267: data = 8'h06;
      17'd14268: data = 8'h0d;
      17'd14269: data = 8'h13;
      17'd14270: data = 8'h16;
      17'd14271: data = 8'h1b;
      17'd14272: data = 8'h1f;
      17'd14273: data = 8'h1f;
      17'd14274: data = 8'h1f;
      17'd14275: data = 8'h1a;
      17'd14276: data = 8'h0e;
      17'd14277: data = 8'h0d;
      17'd14278: data = 8'h09;
      17'd14279: data = 8'h06;
      17'd14280: data = 8'h0d;
      17'd14281: data = 8'h15;
      17'd14282: data = 8'h1a;
      17'd14283: data = 8'h16;
      17'd14284: data = 8'h0a;
      17'd14285: data = 8'h01;
      17'd14286: data = 8'h00;
      17'd14287: data = 8'h00;
      17'd14288: data = 8'hfd;
      17'd14289: data = 8'hfd;
      17'd14290: data = 8'hfd;
      17'd14291: data = 8'hf9;
      17'd14292: data = 8'hf9;
      17'd14293: data = 8'hf2;
      17'd14294: data = 8'hec;
      17'd14295: data = 8'heb;
      17'd14296: data = 8'he7;
      17'd14297: data = 8'heb;
      17'd14298: data = 8'hed;
      17'd14299: data = 8'heb;
      17'd14300: data = 8'hec;
      17'd14301: data = 8'hed;
      17'd14302: data = 8'hef;
      17'd14303: data = 8'hec;
      17'd14304: data = 8'heb;
      17'd14305: data = 8'he4;
      17'd14306: data = 8'hde;
      17'd14307: data = 8'he0;
      17'd14308: data = 8'he3;
      17'd14309: data = 8'he4;
      17'd14310: data = 8'hf1;
      17'd14311: data = 8'h02;
      17'd14312: data = 8'h04;
      17'd14313: data = 8'h00;
      17'd14314: data = 8'hfa;
      17'd14315: data = 8'hf4;
      17'd14316: data = 8'hfd;
      17'd14317: data = 8'hfc;
      17'd14318: data = 8'hf6;
      17'd14319: data = 8'hfd;
      17'd14320: data = 8'h05;
      17'd14321: data = 8'h06;
      17'd14322: data = 8'hfd;
      17'd14323: data = 8'h05;
      17'd14324: data = 8'h0c;
      17'd14325: data = 8'h09;
      17'd14326: data = 8'h16;
      17'd14327: data = 8'h1a;
      17'd14328: data = 8'h12;
      17'd14329: data = 8'h1a;
      17'd14330: data = 8'h1c;
      17'd14331: data = 8'h0e;
      17'd14332: data = 8'h1b;
      17'd14333: data = 8'h1e;
      17'd14334: data = 8'h06;
      17'd14335: data = 8'h0d;
      17'd14336: data = 8'h05;
      17'd14337: data = 8'h05;
      17'd14338: data = 8'h1e;
      17'd14339: data = 8'h16;
      17'd14340: data = 8'h13;
      17'd14341: data = 8'h2b;
      17'd14342: data = 8'h27;
      17'd14343: data = 8'h0c;
      17'd14344: data = 8'h01;
      17'd14345: data = 8'hf5;
      17'd14346: data = 8'hde;
      17'd14347: data = 8'he9;
      17'd14348: data = 8'hfd;
      17'd14349: data = 8'hfe;
      17'd14350: data = 8'h09;
      17'd14351: data = 8'h24;
      17'd14352: data = 8'h1b;
      17'd14353: data = 8'h01;
      17'd14354: data = 8'hfc;
      17'd14355: data = 8'he9;
      17'd14356: data = 8'he3;
      17'd14357: data = 8'hdc;
      17'd14358: data = 8'hda;
      17'd14359: data = 8'hf6;
      17'd14360: data = 8'h01;
      17'd14361: data = 8'h04;
      17'd14362: data = 8'h12;
      17'd14363: data = 8'h0c;
      17'd14364: data = 8'hf5;
      17'd14365: data = 8'hf6;
      17'd14366: data = 8'hfe;
      17'd14367: data = 8'hf5;
      17'd14368: data = 8'hf9;
      17'd14369: data = 8'h05;
      17'd14370: data = 8'h0d;
      17'd14371: data = 8'h06;
      17'd14372: data = 8'h0a;
      17'd14373: data = 8'h11;
      17'd14374: data = 8'hfd;
      17'd14375: data = 8'hf2;
      17'd14376: data = 8'hfd;
      17'd14377: data = 8'h09;
      17'd14378: data = 8'h0c;
      17'd14379: data = 8'h1a;
      17'd14380: data = 8'h26;
      17'd14381: data = 8'h1e;
      17'd14382: data = 8'h16;
      17'd14383: data = 8'h0a;
      17'd14384: data = 8'hfc;
      17'd14385: data = 8'hf2;
      17'd14386: data = 8'hf9;
      17'd14387: data = 8'hfd;
      17'd14388: data = 8'h04;
      17'd14389: data = 8'h0d;
      17'd14390: data = 8'h12;
      17'd14391: data = 8'h1b;
      17'd14392: data = 8'h0d;
      17'd14393: data = 8'hf5;
      17'd14394: data = 8'hf4;
      17'd14395: data = 8'hec;
      17'd14396: data = 8'he3;
      17'd14397: data = 8'hec;
      17'd14398: data = 8'hec;
      17'd14399: data = 8'he9;
      17'd14400: data = 8'hf4;
      17'd14401: data = 8'hf5;
      17'd14402: data = 8'he9;
      17'd14403: data = 8'he4;
      17'd14404: data = 8'he2;
      17'd14405: data = 8'hdc;
      17'd14406: data = 8'hdb;
      17'd14407: data = 8'he2;
      17'd14408: data = 8'he5;
      17'd14409: data = 8'heb;
      17'd14410: data = 8'hec;
      17'd14411: data = 8'he5;
      17'd14412: data = 8'he5;
      17'd14413: data = 8'hdb;
      17'd14414: data = 8'hd8;
      17'd14415: data = 8'he0;
      17'd14416: data = 8'he2;
      17'd14417: data = 8'hec;
      17'd14418: data = 8'hf9;
      17'd14419: data = 8'h00;
      17'd14420: data = 8'h00;
      17'd14421: data = 8'h04;
      17'd14422: data = 8'h00;
      17'd14423: data = 8'hf9;
      17'd14424: data = 8'hfa;
      17'd14425: data = 8'h00;
      17'd14426: data = 8'h09;
      17'd14427: data = 8'h0e;
      17'd14428: data = 8'h16;
      17'd14429: data = 8'h22;
      17'd14430: data = 8'h26;
      17'd14431: data = 8'h23;
      17'd14432: data = 8'h1f;
      17'd14433: data = 8'h1f;
      17'd14434: data = 8'h1a;
      17'd14435: data = 8'h22;
      17'd14436: data = 8'h27;
      17'd14437: data = 8'h26;
      17'd14438: data = 8'h31;
      17'd14439: data = 8'h34;
      17'd14440: data = 8'h31;
      17'd14441: data = 8'h2d;
      17'd14442: data = 8'h29;
      17'd14443: data = 8'h22;
      17'd14444: data = 8'h22;
      17'd14445: data = 8'h23;
      17'd14446: data = 8'h24;
      17'd14447: data = 8'h2c;
      17'd14448: data = 8'h29;
      17'd14449: data = 8'h24;
      17'd14450: data = 8'h22;
      17'd14451: data = 8'h15;
      17'd14452: data = 8'h0d;
      17'd14453: data = 8'h09;
      17'd14454: data = 8'h05;
      17'd14455: data = 8'h05;
      17'd14456: data = 8'h0a;
      17'd14457: data = 8'h09;
      17'd14458: data = 8'h04;
      17'd14459: data = 8'h06;
      17'd14460: data = 8'h00;
      17'd14461: data = 8'hf4;
      17'd14462: data = 8'hed;
      17'd14463: data = 8'he7;
      17'd14464: data = 8'he4;
      17'd14465: data = 8'hec;
      17'd14466: data = 8'hec;
      17'd14467: data = 8'he7;
      17'd14468: data = 8'hec;
      17'd14469: data = 8'heb;
      17'd14470: data = 8'he2;
      17'd14471: data = 8'hdc;
      17'd14472: data = 8'hda;
      17'd14473: data = 8'hdb;
      17'd14474: data = 8'hdc;
      17'd14475: data = 8'hd6;
      17'd14476: data = 8'hdb;
      17'd14477: data = 8'he2;
      17'd14478: data = 8'he2;
      17'd14479: data = 8'hde;
      17'd14480: data = 8'hdc;
      17'd14481: data = 8'hdc;
      17'd14482: data = 8'hd8;
      17'd14483: data = 8'hda;
      17'd14484: data = 8'he0;
      17'd14485: data = 8'he4;
      17'd14486: data = 8'heb;
      17'd14487: data = 8'hed;
      17'd14488: data = 8'hf2;
      17'd14489: data = 8'hf4;
      17'd14490: data = 8'hf5;
      17'd14491: data = 8'hf4;
      17'd14492: data = 8'hf1;
      17'd14493: data = 8'hf4;
      17'd14494: data = 8'hfa;
      17'd14495: data = 8'hfd;
      17'd14496: data = 8'h00;
      17'd14497: data = 8'hfe;
      17'd14498: data = 8'h01;
      17'd14499: data = 8'h02;
      17'd14500: data = 8'h00;
      17'd14501: data = 8'h00;
      17'd14502: data = 8'h05;
      17'd14503: data = 8'h09;
      17'd14504: data = 8'h05;
      17'd14505: data = 8'h09;
      17'd14506: data = 8'h09;
      17'd14507: data = 8'h0a;
      17'd14508: data = 8'h0e;
      17'd14509: data = 8'h0a;
      17'd14510: data = 8'h06;
      17'd14511: data = 8'h05;
      17'd14512: data = 8'h05;
      17'd14513: data = 8'h05;
      17'd14514: data = 8'h02;
      17'd14515: data = 8'h05;
      17'd14516: data = 8'h05;
      17'd14517: data = 8'h05;
      17'd14518: data = 8'h09;
      17'd14519: data = 8'h01;
      17'd14520: data = 8'h00;
      17'd14521: data = 8'hfd;
      17'd14522: data = 8'hf6;
      17'd14523: data = 8'hf6;
      17'd14524: data = 8'hf9;
      17'd14525: data = 8'hfc;
      17'd14526: data = 8'hfd;
      17'd14527: data = 8'hfe;
      17'd14528: data = 8'hfc;
      17'd14529: data = 8'hf9;
      17'd14530: data = 8'hf5;
      17'd14531: data = 8'hf4;
      17'd14532: data = 8'hf5;
      17'd14533: data = 8'hfc;
      17'd14534: data = 8'hf6;
      17'd14535: data = 8'hf2;
      17'd14536: data = 8'hf5;
      17'd14537: data = 8'hf6;
      17'd14538: data = 8'hf4;
      17'd14539: data = 8'hf4;
      17'd14540: data = 8'hf2;
      17'd14541: data = 8'hf1;
      17'd14542: data = 8'hfc;
      17'd14543: data = 8'hfe;
      17'd14544: data = 8'hf6;
      17'd14545: data = 8'hf9;
      17'd14546: data = 8'hf5;
      17'd14547: data = 8'hed;
      17'd14548: data = 8'h05;
      17'd14549: data = 8'h23;
      17'd14550: data = 8'h01;
      17'd14551: data = 8'he7;
      17'd14552: data = 8'hfa;
      17'd14553: data = 8'hfa;
      17'd14554: data = 8'h00;
      17'd14555: data = 8'h1b;
      17'd14556: data = 8'h12;
      17'd14557: data = 8'hf6;
      17'd14558: data = 8'hfe;
      17'd14559: data = 8'h12;
      17'd14560: data = 8'h1c;
      17'd14561: data = 8'h09;
      17'd14562: data = 8'hfd;
      17'd14563: data = 8'h15;
      17'd14564: data = 8'h09;
      17'd14565: data = 8'hfd;
      17'd14566: data = 8'h16;
      17'd14567: data = 8'h11;
      17'd14568: data = 8'h00;
      17'd14569: data = 8'h0d;
      17'd14570: data = 8'h15;
      17'd14571: data = 8'h02;
      17'd14572: data = 8'h09;
      17'd14573: data = 8'h22;
      17'd14574: data = 8'h01;
      17'd14575: data = 8'hfd;
      17'd14576: data = 8'h12;
      17'd14577: data = 8'h0d;
      17'd14578: data = 8'h09;
      17'd14579: data = 8'hef;
      17'd14580: data = 8'hfe;
      17'd14581: data = 8'h13;
      17'd14582: data = 8'hf4;
      17'd14583: data = 8'hf9;
      17'd14584: data = 8'h19;
      17'd14585: data = 8'h15;
      17'd14586: data = 8'hfd;
      17'd14587: data = 8'h00;
      17'd14588: data = 8'h02;
      17'd14589: data = 8'hfd;
      17'd14590: data = 8'hf5;
      17'd14591: data = 8'hed;
      17'd14592: data = 8'hec;
      17'd14593: data = 8'hef;
      17'd14594: data = 8'hfe;
      17'd14595: data = 8'h11;
      17'd14596: data = 8'h01;
      17'd14597: data = 8'hef;
      17'd14598: data = 8'hfc;
      17'd14599: data = 8'h05;
      17'd14600: data = 8'hf6;
      17'd14601: data = 8'hf9;
      17'd14602: data = 8'h0a;
      17'd14603: data = 8'hf9;
      17'd14604: data = 8'hf1;
      17'd14605: data = 8'hfe;
      17'd14606: data = 8'hfd;
      17'd14607: data = 8'hfa;
      17'd14608: data = 8'hfc;
      17'd14609: data = 8'hfe;
      17'd14610: data = 8'hfe;
      17'd14611: data = 8'hfe;
      17'd14612: data = 8'h0e;
      17'd14613: data = 8'h16;
      17'd14614: data = 8'h11;
      17'd14615: data = 8'h0d;
      17'd14616: data = 8'h11;
      17'd14617: data = 8'h04;
      17'd14618: data = 8'hfa;
      17'd14619: data = 8'h01;
      17'd14620: data = 8'h00;
      17'd14621: data = 8'hfd;
      17'd14622: data = 8'h04;
      17'd14623: data = 8'h09;
      17'd14624: data = 8'h0d;
      17'd14625: data = 8'h0d;
      17'd14626: data = 8'h11;
      17'd14627: data = 8'h0c;
      17'd14628: data = 8'hfe;
      17'd14629: data = 8'h09;
      17'd14630: data = 8'h0d;
      17'd14631: data = 8'h02;
      17'd14632: data = 8'h01;
      17'd14633: data = 8'h04;
      17'd14634: data = 8'h01;
      17'd14635: data = 8'hfa;
      17'd14636: data = 8'hfd;
      17'd14637: data = 8'hfd;
      17'd14638: data = 8'hf9;
      17'd14639: data = 8'hfe;
      17'd14640: data = 8'h01;
      17'd14641: data = 8'hfc;
      17'd14642: data = 8'hf9;
      17'd14643: data = 8'hfd;
      17'd14644: data = 8'hfc;
      17'd14645: data = 8'hf1;
      17'd14646: data = 8'hed;
      17'd14647: data = 8'hf2;
      17'd14648: data = 8'hef;
      17'd14649: data = 8'heb;
      17'd14650: data = 8'hf5;
      17'd14651: data = 8'hf6;
      17'd14652: data = 8'hf2;
      17'd14653: data = 8'hf6;
      17'd14654: data = 8'hf6;
      17'd14655: data = 8'hf4;
      17'd14656: data = 8'hf5;
      17'd14657: data = 8'hf9;
      17'd14658: data = 8'hf9;
      17'd14659: data = 8'hf6;
      17'd14660: data = 8'hfc;
      17'd14661: data = 8'h00;
      17'd14662: data = 8'hf9;
      17'd14663: data = 8'hf9;
      17'd14664: data = 8'h00;
      17'd14665: data = 8'h02;
      17'd14666: data = 8'h00;
      17'd14667: data = 8'h02;
      17'd14668: data = 8'h09;
      17'd14669: data = 8'h0a;
      17'd14670: data = 8'h0c;
      17'd14671: data = 8'h0a;
      17'd14672: data = 8'h09;
      17'd14673: data = 8'h09;
      17'd14674: data = 8'h05;
      17'd14675: data = 8'h05;
      17'd14676: data = 8'h0d;
      17'd14677: data = 8'h11;
      17'd14678: data = 8'h0d;
      17'd14679: data = 8'h0a;
      17'd14680: data = 8'h13;
      17'd14681: data = 8'h1c;
      17'd14682: data = 8'h15;
      17'd14683: data = 8'h0c;
      17'd14684: data = 8'h0c;
      17'd14685: data = 8'h12;
      17'd14686: data = 8'h12;
      17'd14687: data = 8'h0e;
      17'd14688: data = 8'h0e;
      17'd14689: data = 8'h0d;
      17'd14690: data = 8'h0c;
      17'd14691: data = 8'h0e;
      17'd14692: data = 8'h11;
      17'd14693: data = 8'h06;
      17'd14694: data = 8'h04;
      17'd14695: data = 8'h06;
      17'd14696: data = 8'h06;
      17'd14697: data = 8'h0e;
      17'd14698: data = 8'h0a;
      17'd14699: data = 8'hfd;
      17'd14700: data = 8'hfa;
      17'd14701: data = 8'h04;
      17'd14702: data = 8'h06;
      17'd14703: data = 8'hfe;
      17'd14704: data = 8'hf6;
      17'd14705: data = 8'hf4;
      17'd14706: data = 8'hfd;
      17'd14707: data = 8'h02;
      17'd14708: data = 8'hfe;
      17'd14709: data = 8'hfc;
      17'd14710: data = 8'hf5;
      17'd14711: data = 8'hf5;
      17'd14712: data = 8'hfa;
      17'd14713: data = 8'hf4;
      17'd14714: data = 8'hf1;
      17'd14715: data = 8'hf5;
      17'd14716: data = 8'hf5;
      17'd14717: data = 8'hf1;
      17'd14718: data = 8'heb;
      17'd14719: data = 8'hed;
      17'd14720: data = 8'hef;
      17'd14721: data = 8'hf6;
      17'd14722: data = 8'h01;
      17'd14723: data = 8'hfa;
      17'd14724: data = 8'he9;
      17'd14725: data = 8'heb;
      17'd14726: data = 8'hf4;
      17'd14727: data = 8'hf5;
      17'd14728: data = 8'hf4;
      17'd14729: data = 8'hed;
      17'd14730: data = 8'he9;
      17'd14731: data = 8'he7;
      17'd14732: data = 8'hf9;
      17'd14733: data = 8'h01;
      17'd14734: data = 8'he0;
      17'd14735: data = 8'he5;
      17'd14736: data = 8'h09;
      17'd14737: data = 8'hf2;
      17'd14738: data = 8'he3;
      17'd14739: data = 8'hfe;
      17'd14740: data = 8'hfa;
      17'd14741: data = 8'he7;
      17'd14742: data = 8'hf2;
      17'd14743: data = 8'hfd;
      17'd14744: data = 8'h02;
      17'd14745: data = 8'hef;
      17'd14746: data = 8'he3;
      17'd14747: data = 8'hfc;
      17'd14748: data = 8'hed;
      17'd14749: data = 8'heb;
      17'd14750: data = 8'h16;
      17'd14751: data = 8'hfe;
      17'd14752: data = 8'he0;
      17'd14753: data = 8'hf9;
      17'd14754: data = 8'h11;
      17'd14755: data = 8'h02;
      17'd14756: data = 8'hd6;
      17'd14757: data = 8'he4;
      17'd14758: data = 8'h19;
      17'd14759: data = 8'h1e;
      17'd14760: data = 8'hf2;
      17'd14761: data = 8'hce;
      17'd14762: data = 8'hfe;
      17'd14763: data = 8'h29;
      17'd14764: data = 8'hfd;
      17'd14765: data = 8'he3;
      17'd14766: data = 8'h01;
      17'd14767: data = 8'h0c;
      17'd14768: data = 8'h05;
      17'd14769: data = 8'hf5;
      17'd14770: data = 8'hdb;
      17'd14771: data = 8'h11;
      17'd14772: data = 8'h43;
      17'd14773: data = 8'he0;
      17'd14774: data = 8'hd5;
      17'd14775: data = 8'h27;
      17'd14776: data = 8'hf4;
      17'd14777: data = 8'h1b;
      17'd14778: data = 8'heb;
      17'd14779: data = 8'hc1;
      17'd14780: data = 8'h63;
      17'd14781: data = 8'h22;
      17'd14782: data = 8'ha4;
      17'd14783: data = 8'h02;
      17'd14784: data = 8'h2c;
      17'd14785: data = 8'hf6;
      17'd14786: data = 8'hf5;
      17'd14787: data = 8'h13;
      17'd14788: data = 8'hec;
      17'd14789: data = 8'hf9;
      17'd14790: data = 8'h24;
      17'd14791: data = 8'he9;
      17'd14792: data = 8'h0c;
      17'd14793: data = 8'h12;
      17'd14794: data = 8'hd8;
      17'd14795: data = 8'h1e;
      17'd14796: data = 8'h0d;
      17'd14797: data = 8'he7;
      17'd14798: data = 8'h1c;
      17'd14799: data = 8'hf9;
      17'd14800: data = 8'he3;
      17'd14801: data = 8'h24;
      17'd14802: data = 8'hfa;
      17'd14803: data = 8'h13;
      17'd14804: data = 8'h11;
      17'd14805: data = 8'hb3;
      17'd14806: data = 8'h29;
      17'd14807: data = 8'h31;
      17'd14808: data = 8'hd3;
      17'd14809: data = 8'h13;
      17'd14810: data = 8'hf6;
      17'd14811: data = 8'h22;
      17'd14812: data = 8'h09;
      17'd14813: data = 8'hc1;
      17'd14814: data = 8'h42;
      17'd14815: data = 8'h0a;
      17'd14816: data = 8'hc5;
      17'd14817: data = 8'h3d;
      17'd14818: data = 8'h00;
      17'd14819: data = 8'hd5;
      17'd14820: data = 8'h35;
      17'd14821: data = 8'hf1;
      17'd14822: data = 8'hfa;
      17'd14823: data = 8'h1e;
      17'd14824: data = 8'he2;
      17'd14825: data = 8'h09;
      17'd14826: data = 8'h1c;
      17'd14827: data = 8'hf1;
      17'd14828: data = 8'hfe;
      17'd14829: data = 8'h11;
      17'd14830: data = 8'hf1;
      17'd14831: data = 8'h04;
      17'd14832: data = 8'h12;
      17'd14833: data = 8'he5;
      17'd14834: data = 8'h12;
      17'd14835: data = 8'h12;
      17'd14836: data = 8'hdc;
      17'd14837: data = 8'h15;
      17'd14838: data = 8'h19;
      17'd14839: data = 8'hdc;
      17'd14840: data = 8'h16;
      17'd14841: data = 8'h13;
      17'd14842: data = 8'hdc;
      17'd14843: data = 8'h1c;
      17'd14844: data = 8'h11;
      17'd14845: data = 8'hd3;
      17'd14846: data = 8'h16;
      17'd14847: data = 8'h0d;
      17'd14848: data = 8'hed;
      17'd14849: data = 8'h0c;
      17'd14850: data = 8'h09;
      17'd14851: data = 8'hf1;
      17'd14852: data = 8'h00;
      17'd14853: data = 8'h11;
      17'd14854: data = 8'hf5;
      17'd14855: data = 8'h02;
      17'd14856: data = 8'h0c;
      17'd14857: data = 8'hfc;
      17'd14858: data = 8'hfe;
      17'd14859: data = 8'hfa;
      17'd14860: data = 8'h11;
      17'd14861: data = 8'h0e;
      17'd14862: data = 8'hdb;
      17'd14863: data = 8'h0c;
      17'd14864: data = 8'h1f;
      17'd14865: data = 8'hdb;
      17'd14866: data = 8'h09;
      17'd14867: data = 8'h1a;
      17'd14868: data = 8'he3;
      17'd14869: data = 8'h06;
      17'd14870: data = 8'h11;
      17'd14871: data = 8'hec;
      17'd14872: data = 8'h02;
      17'd14873: data = 8'h0c;
      17'd14874: data = 8'hfe;
      17'd14875: data = 8'h0e;
      17'd14876: data = 8'hf9;
      17'd14877: data = 8'hf2;
      17'd14878: data = 8'h19;
      17'd14879: data = 8'h05;
      17'd14880: data = 8'hf9;
      17'd14881: data = 8'h0a;
      17'd14882: data = 8'h06;
      17'd14883: data = 8'h00;
      17'd14884: data = 8'h02;
      17'd14885: data = 8'h0e;
      17'd14886: data = 8'h09;
      17'd14887: data = 8'hfc;
      17'd14888: data = 8'h01;
      17'd14889: data = 8'h09;
      17'd14890: data = 8'h09;
      17'd14891: data = 8'h04;
      17'd14892: data = 8'hfd;
      17'd14893: data = 8'h05;
      17'd14894: data = 8'h02;
      17'd14895: data = 8'h04;
      17'd14896: data = 8'h06;
      17'd14897: data = 8'hfe;
      17'd14898: data = 8'h01;
      17'd14899: data = 8'h05;
      17'd14900: data = 8'hfd;
      17'd14901: data = 8'h02;
      17'd14902: data = 8'h04;
      17'd14903: data = 8'hf5;
      17'd14904: data = 8'h02;
      17'd14905: data = 8'h05;
      17'd14906: data = 8'hfc;
      17'd14907: data = 8'hfe;
      17'd14908: data = 8'hfa;
      17'd14909: data = 8'hf1;
      17'd14910: data = 8'h00;
      17'd14911: data = 8'h04;
      17'd14912: data = 8'hf6;
      17'd14913: data = 8'hf5;
      17'd14914: data = 8'hf5;
      17'd14915: data = 8'hfc;
      17'd14916: data = 8'h01;
      17'd14917: data = 8'hf1;
      17'd14918: data = 8'hf2;
      17'd14919: data = 8'h06;
      17'd14920: data = 8'hfe;
      17'd14921: data = 8'hf5;
      17'd14922: data = 8'hf4;
      17'd14923: data = 8'hf4;
      17'd14924: data = 8'h09;
      17'd14925: data = 8'hf6;
      17'd14926: data = 8'hed;
      17'd14927: data = 8'h09;
      17'd14928: data = 8'hed;
      17'd14929: data = 8'he5;
      17'd14930: data = 8'h0c;
      17'd14931: data = 8'hfe;
      17'd14932: data = 8'hfc;
      17'd14933: data = 8'h00;
      17'd14934: data = 8'he4;
      17'd14935: data = 8'hfe;
      17'd14936: data = 8'h11;
      17'd14937: data = 8'hf6;
      17'd14938: data = 8'hfc;
      17'd14939: data = 8'hfe;
      17'd14940: data = 8'hec;
      17'd14941: data = 8'h06;
      17'd14942: data = 8'h11;
      17'd14943: data = 8'hf1;
      17'd14944: data = 8'h09;
      17'd14945: data = 8'hfc;
      17'd14946: data = 8'hf6;
      17'd14947: data = 8'h16;
      17'd14948: data = 8'hfd;
      17'd14949: data = 8'hfe;
      17'd14950: data = 8'h15;
      17'd14951: data = 8'hec;
      17'd14952: data = 8'hfa;
      17'd14953: data = 8'h24;
      17'd14954: data = 8'hf6;
      17'd14955: data = 8'hf6;
      17'd14956: data = 8'h09;
      17'd14957: data = 8'hf5;
      17'd14958: data = 8'h09;
      17'd14959: data = 8'h0d;
      17'd14960: data = 8'hf9;
      17'd14961: data = 8'h01;
      17'd14962: data = 8'h02;
      17'd14963: data = 8'hfa;
      17'd14964: data = 8'hfe;
      17'd14965: data = 8'h05;
      17'd14966: data = 8'h05;
      17'd14967: data = 8'hfc;
      17'd14968: data = 8'hf4;
      17'd14969: data = 8'hfc;
      17'd14970: data = 8'h05;
      17'd14971: data = 8'hfd;
      17'd14972: data = 8'hf6;
      17'd14973: data = 8'h00;
      17'd14974: data = 8'hed;
      17'd14975: data = 8'hed;
      17'd14976: data = 8'h12;
      17'd14977: data = 8'h02;
      17'd14978: data = 8'hdb;
      17'd14979: data = 8'h05;
      17'd14980: data = 8'h09;
      17'd14981: data = 8'hda;
      17'd14982: data = 8'h09;
      17'd14983: data = 8'h0d;
      17'd14984: data = 8'he3;
      17'd14985: data = 8'hfc;
      17'd14986: data = 8'hfa;
      17'd14987: data = 8'hfa;
      17'd14988: data = 8'h0a;
      17'd14989: data = 8'he3;
      17'd14990: data = 8'hfa;
      17'd14991: data = 8'h15;
      17'd14992: data = 8'hda;
      17'd14993: data = 8'hfc;
      17'd14994: data = 8'h24;
      17'd14995: data = 8'he2;
      17'd14996: data = 8'he5;
      17'd14997: data = 8'h12;
      17'd14998: data = 8'hfd;
      17'd14999: data = 8'hf4;
      17'd15000: data = 8'h01;
      17'd15001: data = 8'h09;
      17'd15002: data = 8'hf9;
      17'd15003: data = 8'he7;
      17'd15004: data = 8'h06;
      17'd15005: data = 8'h09;
      17'd15006: data = 8'hf9;
      17'd15007: data = 8'h11;
      17'd15008: data = 8'hf6;
      17'd15009: data = 8'he5;
      17'd15010: data = 8'h13;
      17'd15011: data = 8'h11;
      17'd15012: data = 8'hed;
      17'd15013: data = 8'hfd;
      17'd15014: data = 8'h12;
      17'd15015: data = 8'hef;
      17'd15016: data = 8'hf6;
      17'd15017: data = 8'h1e;
      17'd15018: data = 8'hf6;
      17'd15019: data = 8'hf6;
      17'd15020: data = 8'h05;
      17'd15021: data = 8'hed;
      17'd15022: data = 8'h13;
      17'd15023: data = 8'h0e;
      17'd15024: data = 8'hde;
      17'd15025: data = 8'h06;
      17'd15026: data = 8'h0e;
      17'd15027: data = 8'he9;
      17'd15028: data = 8'h06;
      17'd15029: data = 8'h04;
      17'd15030: data = 8'hed;
      17'd15031: data = 8'h0e;
      17'd15032: data = 8'hfa;
      17'd15033: data = 8'he3;
      17'd15034: data = 8'h11;
      17'd15035: data = 8'h00;
      17'd15036: data = 8'heb;
      17'd15037: data = 8'h0a;
      17'd15038: data = 8'h04;
      17'd15039: data = 8'he9;
      17'd15040: data = 8'h02;
      17'd15041: data = 8'h0c;
      17'd15042: data = 8'hed;
      17'd15043: data = 8'hfa;
      17'd15044: data = 8'h06;
      17'd15045: data = 8'hfd;
      17'd15046: data = 8'hf6;
      17'd15047: data = 8'hfc;
      17'd15048: data = 8'hf4;
      17'd15049: data = 8'hfc;
      17'd15050: data = 8'h0d;
      17'd15051: data = 8'h00;
      17'd15052: data = 8'he4;
      17'd15053: data = 8'hf9;
      17'd15054: data = 8'h1c;
      17'd15055: data = 8'hfd;
      17'd15056: data = 8'he4;
      17'd15057: data = 8'h02;
      17'd15058: data = 8'hfe;
      17'd15059: data = 8'hf9;
      17'd15060: data = 8'h1e;
      17'd15061: data = 8'hfc;
      17'd15062: data = 8'hdb;
      17'd15063: data = 8'hfd;
      17'd15064: data = 8'h0e;
      17'd15065: data = 8'h0d;
      17'd15066: data = 8'h0e;
      17'd15067: data = 8'hf4;
      17'd15068: data = 8'hde;
      17'd15069: data = 8'h04;
      17'd15070: data = 8'h1f;
      17'd15071: data = 8'h04;
      17'd15072: data = 8'h04;
      17'd15073: data = 8'hf2;
      17'd15074: data = 8'hde;
      17'd15075: data = 8'h1f;
      17'd15076: data = 8'h23;
      17'd15077: data = 8'he5;
      17'd15078: data = 8'hec;
      17'd15079: data = 8'h1e;
      17'd15080: data = 8'hed;
      17'd15081: data = 8'h01;
      17'd15082: data = 8'h24;
      17'd15083: data = 8'hce;
      17'd15084: data = 8'h05;
      17'd15085: data = 8'h33;
      17'd15086: data = 8'hd1;
      17'd15087: data = 8'h01;
      17'd15088: data = 8'h29;
      17'd15089: data = 8'hdb;
      17'd15090: data = 8'h02;
      17'd15091: data = 8'h15;
      17'd15092: data = 8'he3;
      17'd15093: data = 8'h01;
      17'd15094: data = 8'h0d;
      17'd15095: data = 8'hfc;
      17'd15096: data = 8'h09;
      17'd15097: data = 8'hf4;
      17'd15098: data = 8'hfe;
      17'd15099: data = 8'h13;
      17'd15100: data = 8'hf4;
      17'd15101: data = 8'h09;
      17'd15102: data = 8'h02;
      17'd15103: data = 8'h02;
      17'd15104: data = 8'h09;
      17'd15105: data = 8'hf4;
      17'd15106: data = 8'h19;
      17'd15107: data = 8'h0c;
      17'd15108: data = 8'hed;
      17'd15109: data = 8'h1b;
      17'd15110: data = 8'h04;
      17'd15111: data = 8'he0;
      17'd15112: data = 8'h35;
      17'd15113: data = 8'h11;
      17'd15114: data = 8'hce;
      17'd15115: data = 8'h36;
      17'd15116: data = 8'h05;
      17'd15117: data = 8'hd5;
      17'd15118: data = 8'h4e;
      17'd15119: data = 8'h09;
      17'd15120: data = 8'hc9;
      17'd15121: data = 8'h26;
      17'd15122: data = 8'h1b;
      17'd15123: data = 8'hfd;
      17'd15124: data = 8'h0e;
      17'd15125: data = 8'h13;
      17'd15126: data = 8'hfd;
      17'd15127: data = 8'hf1;
      17'd15128: data = 8'h26;
      17'd15129: data = 8'h24;
      17'd15130: data = 8'hda;
      17'd15131: data = 8'hf9;
      17'd15132: data = 8'h2b;
      17'd15133: data = 8'hf2;
      17'd15134: data = 8'h02;
      17'd15135: data = 8'h16;
      17'd15136: data = 8'hf2;
      17'd15137: data = 8'hfd;
      17'd15138: data = 8'hfd;
      17'd15139: data = 8'h1a;
      17'd15140: data = 8'h0e;
      17'd15141: data = 8'hd2;
      17'd15142: data = 8'h12;
      17'd15143: data = 8'h1c;
      17'd15144: data = 8'hd3;
      17'd15145: data = 8'h0d;
      17'd15146: data = 8'h0e;
      17'd15147: data = 8'hed;
      17'd15148: data = 8'h0c;
      17'd15149: data = 8'he9;
      17'd15150: data = 8'hf5;
      17'd15151: data = 8'h0e;
      17'd15152: data = 8'hfa;
      17'd15153: data = 8'hf9;
      17'd15154: data = 8'h0e;
      17'd15155: data = 8'hf4;
      17'd15156: data = 8'hd8;
      17'd15157: data = 8'h16;
      17'd15158: data = 8'h13;
      17'd15159: data = 8'hef;
      17'd15160: data = 8'h05;
      17'd15161: data = 8'hef;
      17'd15162: data = 8'he3;
      17'd15163: data = 8'h22;
      17'd15164: data = 8'h15;
      17'd15165: data = 8'he5;
      17'd15166: data = 8'hf4;
      17'd15167: data = 8'h0d;
      17'd15168: data = 8'h09;
      17'd15169: data = 8'hfd;
      17'd15170: data = 8'hf6;
      17'd15171: data = 8'h16;
      17'd15172: data = 8'h0e;
      17'd15173: data = 8'hda;
      17'd15174: data = 8'h0d;
      17'd15175: data = 8'h1f;
      17'd15176: data = 8'hfa;
      17'd15177: data = 8'hfc;
      17'd15178: data = 8'h05;
      17'd15179: data = 8'h09;
      17'd15180: data = 8'hf4;
      17'd15181: data = 8'h06;
      17'd15182: data = 8'h29;
      17'd15183: data = 8'hf6;
      17'd15184: data = 8'hdb;
      17'd15185: data = 8'h16;
      17'd15186: data = 8'h15;
      17'd15187: data = 8'he9;
      17'd15188: data = 8'h11;
      17'd15189: data = 8'h1c;
      17'd15190: data = 8'hce;
      17'd15191: data = 8'hf6;
      17'd15192: data = 8'h34;
      17'd15193: data = 8'hf5;
      17'd15194: data = 8'hd8;
      17'd15195: data = 8'h01;
      17'd15196: data = 8'h22;
      17'd15197: data = 8'hf2;
      17'd15198: data = 8'hda;
      17'd15199: data = 8'h0d;
      17'd15200: data = 8'h0e;
      17'd15201: data = 8'hf2;
      17'd15202: data = 8'hf5;
      17'd15203: data = 8'hef;
      17'd15204: data = 8'hf6;
      17'd15205: data = 8'h11;
      17'd15206: data = 8'hf2;
      17'd15207: data = 8'he7;
      17'd15208: data = 8'hfe;
      17'd15209: data = 8'hec;
      17'd15210: data = 8'hf9;
      17'd15211: data = 8'h0d;
      17'd15212: data = 8'he4;
      17'd15213: data = 8'hf4;
      17'd15214: data = 8'h13;
      17'd15215: data = 8'hd3;
      17'd15216: data = 8'hde;
      17'd15217: data = 8'h33;
      17'd15218: data = 8'hf9;
      17'd15219: data = 8'hc1;
      17'd15220: data = 8'h11;
      17'd15221: data = 8'h0e;
      17'd15222: data = 8'hce;
      17'd15223: data = 8'h0a;
      17'd15224: data = 8'h06;
      17'd15225: data = 8'hd1;
      17'd15226: data = 8'h09;
      17'd15227: data = 8'h15;
      17'd15228: data = 8'hd6;
      17'd15229: data = 8'hf5;
      17'd15230: data = 8'h13;
      17'd15231: data = 8'hec;
      17'd15232: data = 8'hf5;
      17'd15233: data = 8'h05;
      17'd15234: data = 8'hec;
      17'd15235: data = 8'h0c;
      17'd15236: data = 8'h09;
      17'd15237: data = 8'hda;
      17'd15238: data = 8'h06;
      17'd15239: data = 8'h0d;
      17'd15240: data = 8'hec;
      17'd15241: data = 8'h05;
      17'd15242: data = 8'h09;
      17'd15243: data = 8'hed;
      17'd15244: data = 8'h09;
      17'd15245: data = 8'h06;
      17'd15246: data = 8'he4;
      17'd15247: data = 8'h09;
      17'd15248: data = 8'h1a;
      17'd15249: data = 8'hf6;
      17'd15250: data = 8'he9;
      17'd15251: data = 8'h11;
      17'd15252: data = 8'h0a;
      17'd15253: data = 8'heb;
      17'd15254: data = 8'hfd;
      17'd15255: data = 8'h04;
      17'd15256: data = 8'h06;
      17'd15257: data = 8'h04;
      17'd15258: data = 8'hec;
      17'd15259: data = 8'hf5;
      17'd15260: data = 8'h0a;
      17'd15261: data = 8'h11;
      17'd15262: data = 8'h05;
      17'd15263: data = 8'he0;
      17'd15264: data = 8'heb;
      17'd15265: data = 8'h24;
      17'd15266: data = 8'h1a;
      17'd15267: data = 8'hd6;
      17'd15268: data = 8'hf2;
      17'd15269: data = 8'h0a;
      17'd15270: data = 8'h04;
      17'd15271: data = 8'h0e;
      17'd15272: data = 8'hef;
      17'd15273: data = 8'hec;
      17'd15274: data = 8'h04;
      17'd15275: data = 8'h04;
      17'd15276: data = 8'h00;
      17'd15277: data = 8'h0a;
      17'd15278: data = 8'heb;
      17'd15279: data = 8'hec;
      17'd15280: data = 8'h1a;
      17'd15281: data = 8'hfd;
      17'd15282: data = 8'hdb;
      17'd15283: data = 8'h1f;
      17'd15284: data = 8'h0c;
      17'd15285: data = 8'hb9;
      17'd15286: data = 8'h11;
      17'd15287: data = 8'h2d;
      17'd15288: data = 8'he4;
      17'd15289: data = 8'heb;
      17'd15290: data = 8'h06;
      17'd15291: data = 8'h00;
      17'd15292: data = 8'hf6;
      17'd15293: data = 8'hfe;
      17'd15294: data = 8'h01;
      17'd15295: data = 8'h02;
      17'd15296: data = 8'hf9;
      17'd15297: data = 8'heb;
      17'd15298: data = 8'h0a;
      17'd15299: data = 8'h11;
      17'd15300: data = 8'hec;
      17'd15301: data = 8'hfa;
      17'd15302: data = 8'hfd;
      17'd15303: data = 8'hfc;
      17'd15304: data = 8'h16;
      17'd15305: data = 8'h02;
      17'd15306: data = 8'hdc;
      17'd15307: data = 8'hf9;
      17'd15308: data = 8'h1b;
      17'd15309: data = 8'hf5;
      17'd15310: data = 8'hf1;
      17'd15311: data = 8'h06;
      17'd15312: data = 8'h01;
      17'd15313: data = 8'hf4;
      17'd15314: data = 8'hfd;
      17'd15315: data = 8'h15;
      17'd15316: data = 8'hfe;
      17'd15317: data = 8'he7;
      17'd15318: data = 8'h02;
      17'd15319: data = 8'h0c;
      17'd15320: data = 8'h02;
      17'd15321: data = 8'h02;
      17'd15322: data = 8'hef;
      17'd15323: data = 8'hfc;
      17'd15324: data = 8'h02;
      17'd15325: data = 8'h0d;
      17'd15326: data = 8'hfe;
      17'd15327: data = 8'he9;
      17'd15328: data = 8'h0e;
      17'd15329: data = 8'h15;
      17'd15330: data = 8'he0;
      17'd15331: data = 8'hf9;
      17'd15332: data = 8'h29;
      17'd15333: data = 8'hfa;
      17'd15334: data = 8'he9;
      17'd15335: data = 8'h06;
      17'd15336: data = 8'h0d;
      17'd15337: data = 8'h00;
      17'd15338: data = 8'h02;
      17'd15339: data = 8'hfd;
      17'd15340: data = 8'h02;
      17'd15341: data = 8'h01;
      17'd15342: data = 8'h04;
      17'd15343: data = 8'h1b;
      17'd15344: data = 8'hfd;
      17'd15345: data = 8'heb;
      17'd15346: data = 8'h04;
      17'd15347: data = 8'h23;
      17'd15348: data = 8'h06;
      17'd15349: data = 8'hf4;
      17'd15350: data = 8'h04;
      17'd15351: data = 8'hfc;
      17'd15352: data = 8'h00;
      17'd15353: data = 8'h1f;
      17'd15354: data = 8'h0a;
      17'd15355: data = 8'he4;
      17'd15356: data = 8'h05;
      17'd15357: data = 8'h1a;
      17'd15358: data = 8'h01;
      17'd15359: data = 8'hf1;
      17'd15360: data = 8'h13;
      17'd15361: data = 8'h11;
      17'd15362: data = 8'hde;
      17'd15363: data = 8'h0a;
      17'd15364: data = 8'h22;
      17'd15365: data = 8'heb;
      17'd15366: data = 8'hef;
      17'd15367: data = 8'h19;
      17'd15368: data = 8'h0d;
      17'd15369: data = 8'hec;
      17'd15370: data = 8'hf6;
      17'd15371: data = 8'h13;
      17'd15372: data = 8'h06;
      17'd15373: data = 8'hf6;
      17'd15374: data = 8'h0a;
      17'd15375: data = 8'h05;
      17'd15376: data = 8'he9;
      17'd15377: data = 8'hfd;
      17'd15378: data = 8'h23;
      17'd15379: data = 8'h04;
      17'd15380: data = 8'he0;
      17'd15381: data = 8'h04;
      17'd15382: data = 8'h1a;
      17'd15383: data = 8'hfd;
      17'd15384: data = 8'hf1;
      17'd15385: data = 8'h11;
      17'd15386: data = 8'h0e;
      17'd15387: data = 8'heb;
      17'd15388: data = 8'h04;
      17'd15389: data = 8'h27;
      17'd15390: data = 8'hfa;
      17'd15391: data = 8'he3;
      17'd15392: data = 8'h13;
      17'd15393: data = 8'h19;
      17'd15394: data = 8'hec;
      17'd15395: data = 8'h05;
      17'd15396: data = 8'h19;
      17'd15397: data = 8'hf5;
      17'd15398: data = 8'hfc;
      17'd15399: data = 8'h11;
      17'd15400: data = 8'h12;
      17'd15401: data = 8'hfc;
      17'd15402: data = 8'hf4;
      17'd15403: data = 8'h16;
      17'd15404: data = 8'h19;
      17'd15405: data = 8'hed;
      17'd15406: data = 8'h04;
      17'd15407: data = 8'h15;
      17'd15408: data = 8'hf9;
      17'd15409: data = 8'h0c;
      17'd15410: data = 8'h11;
      17'd15411: data = 8'heb;
      17'd15412: data = 8'h00;
      17'd15413: data = 8'h1e;
      17'd15414: data = 8'h00;
      17'd15415: data = 8'hf5;
      17'd15416: data = 8'hfd;
      17'd15417: data = 8'h0c;
      17'd15418: data = 8'h09;
      17'd15419: data = 8'hfa;
      17'd15420: data = 8'h06;
      17'd15421: data = 8'h09;
      17'd15422: data = 8'heb;
      17'd15423: data = 8'h01;
      17'd15424: data = 8'h16;
      17'd15425: data = 8'hf2;
      17'd15426: data = 8'hf4;
      17'd15427: data = 8'h05;
      17'd15428: data = 8'h11;
      17'd15429: data = 8'he9;
      17'd15430: data = 8'he7;
      17'd15431: data = 8'h22;
      17'd15432: data = 8'hfd;
      17'd15433: data = 8'he7;
      17'd15434: data = 8'hfe;
      17'd15435: data = 8'hf9;
      17'd15436: data = 8'h01;
      17'd15437: data = 8'h02;
      17'd15438: data = 8'hed;
      17'd15439: data = 8'hef;
      17'd15440: data = 8'h09;
      17'd15441: data = 8'h09;
      17'd15442: data = 8'he4;
      17'd15443: data = 8'hf2;
      17'd15444: data = 8'h11;
      17'd15445: data = 8'hf5;
      17'd15446: data = 8'hf2;
      17'd15447: data = 8'h06;
      17'd15448: data = 8'hf4;
      17'd15449: data = 8'hf5;
      17'd15450: data = 8'h0c;
      17'd15451: data = 8'hec;
      17'd15452: data = 8'he9;
      17'd15453: data = 8'h12;
      17'd15454: data = 8'h01;
      17'd15455: data = 8'hec;
      17'd15456: data = 8'hf2;
      17'd15457: data = 8'hfa;
      17'd15458: data = 8'h0c;
      17'd15459: data = 8'hfc;
      17'd15460: data = 8'he5;
      17'd15461: data = 8'h06;
      17'd15462: data = 8'h06;
      17'd15463: data = 8'hfa;
      17'd15464: data = 8'h00;
      17'd15465: data = 8'he7;
      17'd15466: data = 8'h00;
      17'd15467: data = 8'h15;
      17'd15468: data = 8'heb;
      17'd15469: data = 8'hf5;
      17'd15470: data = 8'h13;
      17'd15471: data = 8'hf4;
      17'd15472: data = 8'hfc;
      17'd15473: data = 8'h09;
      17'd15474: data = 8'hf4;
      17'd15475: data = 8'h05;
      17'd15476: data = 8'hfd;
      17'd15477: data = 8'hf6;
      17'd15478: data = 8'h00;
      17'd15479: data = 8'h02;
      17'd15480: data = 8'h12;
      17'd15481: data = 8'hed;
      17'd15482: data = 8'he2;
      17'd15483: data = 8'h13;
      17'd15484: data = 8'h02;
      17'd15485: data = 8'hf1;
      17'd15486: data = 8'h05;
      17'd15487: data = 8'h00;
      17'd15488: data = 8'hfa;
      17'd15489: data = 8'h02;
      17'd15490: data = 8'hfa;
      17'd15491: data = 8'hf1;
      17'd15492: data = 8'h11;
      17'd15493: data = 8'h12;
      17'd15494: data = 8'he5;
      17'd15495: data = 8'hec;
      17'd15496: data = 8'h09;
      17'd15497: data = 8'h0a;
      17'd15498: data = 8'hfe;
      17'd15499: data = 8'hf2;
      17'd15500: data = 8'hf4;
      17'd15501: data = 8'h04;
      17'd15502: data = 8'h02;
      17'd15503: data = 8'hf1;
      17'd15504: data = 8'h05;
      17'd15505: data = 8'h05;
      17'd15506: data = 8'he7;
      17'd15507: data = 8'hf6;
      17'd15508: data = 8'h15;
      17'd15509: data = 8'h0a;
      17'd15510: data = 8'he7;
      17'd15511: data = 8'he9;
      17'd15512: data = 8'hfa;
      17'd15513: data = 8'h11;
      17'd15514: data = 8'h0a;
      17'd15515: data = 8'hec;
      17'd15516: data = 8'hf2;
      17'd15517: data = 8'hfe;
      17'd15518: data = 8'hfa;
      17'd15519: data = 8'h06;
      17'd15520: data = 8'h09;
      17'd15521: data = 8'he3;
      17'd15522: data = 8'hf5;
      17'd15523: data = 8'h1b;
      17'd15524: data = 8'hfa;
      17'd15525: data = 8'hed;
      17'd15526: data = 8'h09;
      17'd15527: data = 8'hf5;
      17'd15528: data = 8'hf1;
      17'd15529: data = 8'h0d;
      17'd15530: data = 8'h00;
      17'd15531: data = 8'he5;
      17'd15532: data = 8'h04;
      17'd15533: data = 8'h0c;
      17'd15534: data = 8'hed;
      17'd15535: data = 8'hfd;
      17'd15536: data = 8'h01;
      17'd15537: data = 8'hf5;
      17'd15538: data = 8'hfc;
      17'd15539: data = 8'h01;
      17'd15540: data = 8'h00;
      17'd15541: data = 8'hfc;
      17'd15542: data = 8'hf1;
      17'd15543: data = 8'h02;
      17'd15544: data = 8'hfe;
      17'd15545: data = 8'hf6;
      17'd15546: data = 8'hfe;
      17'd15547: data = 8'hf1;
      17'd15548: data = 8'h05;
      17'd15549: data = 8'h0d;
      17'd15550: data = 8'hf2;
      17'd15551: data = 8'hf4;
      17'd15552: data = 8'h00;
      17'd15553: data = 8'hfc;
      17'd15554: data = 8'h05;
      17'd15555: data = 8'h16;
      17'd15556: data = 8'hf4;
      17'd15557: data = 8'hd6;
      17'd15558: data = 8'h0a;
      17'd15559: data = 8'h1e;
      17'd15560: data = 8'hf1;
      17'd15561: data = 8'hf6;
      17'd15562: data = 8'h00;
      17'd15563: data = 8'hf2;
      17'd15564: data = 8'h0d;
      17'd15565: data = 8'h0d;
      17'd15566: data = 8'hf2;
      17'd15567: data = 8'h04;
      17'd15568: data = 8'h02;
      17'd15569: data = 8'hf2;
      17'd15570: data = 8'h0c;
      17'd15571: data = 8'h19;
      17'd15572: data = 8'h01;
      17'd15573: data = 8'hf2;
      17'd15574: data = 8'heb;
      17'd15575: data = 8'h0d;
      17'd15576: data = 8'h24;
      17'd15577: data = 8'hf9;
      17'd15578: data = 8'he7;
      17'd15579: data = 8'h05;
      17'd15580: data = 8'h0e;
      17'd15581: data = 8'hfa;
      17'd15582: data = 8'hfa;
      17'd15583: data = 8'h00;
      17'd15584: data = 8'h0c;
      17'd15585: data = 8'h02;
      17'd15586: data = 8'hf5;
      17'd15587: data = 8'h04;
      17'd15588: data = 8'h05;
      17'd15589: data = 8'h00;
      17'd15590: data = 8'h02;
      17'd15591: data = 8'h02;
      17'd15592: data = 8'hfa;
      17'd15593: data = 8'hfd;
      17'd15594: data = 8'h09;
      17'd15595: data = 8'h0d;
      17'd15596: data = 8'hf9;
      17'd15597: data = 8'hec;
      17'd15598: data = 8'hfd;
      17'd15599: data = 8'h12;
      17'd15600: data = 8'h0e;
      17'd15601: data = 8'hf6;
      17'd15602: data = 8'heb;
      17'd15603: data = 8'h0e;
      17'd15604: data = 8'h0d;
      17'd15605: data = 8'hf2;
      17'd15606: data = 8'h11;
      17'd15607: data = 8'h02;
      17'd15608: data = 8'hf1;
      17'd15609: data = 8'h06;
      17'd15610: data = 8'h05;
      17'd15611: data = 8'hfe;
      17'd15612: data = 8'h00;
      17'd15613: data = 8'h00;
      17'd15614: data = 8'h05;
      17'd15615: data = 8'h06;
      17'd15616: data = 8'hfe;
      17'd15617: data = 8'h09;
      17'd15618: data = 8'h05;
      17'd15619: data = 8'h05;
      17'd15620: data = 8'h0a;
      17'd15621: data = 8'h01;
      17'd15622: data = 8'hfe;
      17'd15623: data = 8'h0c;
      17'd15624: data = 8'h0d;
      17'd15625: data = 8'hfd;
      17'd15626: data = 8'hf9;
      17'd15627: data = 8'h0e;
      17'd15628: data = 8'h0a;
      17'd15629: data = 8'h00;
      17'd15630: data = 8'h0d;
      17'd15631: data = 8'h09;
      17'd15632: data = 8'h01;
      17'd15633: data = 8'h09;
      17'd15634: data = 8'h0d;
      17'd15635: data = 8'h09;
      17'd15636: data = 8'h0a;
      17'd15637: data = 8'hf6;
      17'd15638: data = 8'h09;
      17'd15639: data = 8'h16;
      17'd15640: data = 8'hfd;
      17'd15641: data = 8'h09;
      17'd15642: data = 8'h00;
      17'd15643: data = 8'hef;
      17'd15644: data = 8'h19;
      17'd15645: data = 8'h23;
      17'd15646: data = 8'hf1;
      17'd15647: data = 8'hef;
      17'd15648: data = 8'h0e;
      17'd15649: data = 8'h11;
      17'd15650: data = 8'h00;
      17'd15651: data = 8'hf9;
      17'd15652: data = 8'h04;
      17'd15653: data = 8'h00;
      17'd15654: data = 8'hfa;
      17'd15655: data = 8'h05;
      17'd15656: data = 8'h02;
      17'd15657: data = 8'hf6;
      17'd15658: data = 8'h02;
      17'd15659: data = 8'h01;
      17'd15660: data = 8'hef;
      17'd15661: data = 8'h04;
      17'd15662: data = 8'h0e;
      17'd15663: data = 8'hf2;
      17'd15664: data = 8'heb;
      17'd15665: data = 8'h0d;
      17'd15666: data = 8'h06;
      17'd15667: data = 8'hec;
      17'd15668: data = 8'hfc;
      17'd15669: data = 8'h02;
      17'd15670: data = 8'hf6;
      17'd15671: data = 8'hf9;
      17'd15672: data = 8'hfc;
      17'd15673: data = 8'hfd;
      17'd15674: data = 8'h06;
      17'd15675: data = 8'hfa;
      17'd15676: data = 8'hf4;
      17'd15677: data = 8'hfa;
      17'd15678: data = 8'hf1;
      17'd15679: data = 8'h11;
      17'd15680: data = 8'h12;
      17'd15681: data = 8'he4;
      17'd15682: data = 8'hf2;
      17'd15683: data = 8'hfa;
      17'd15684: data = 8'hfa;
      17'd15685: data = 8'h1f;
      17'd15686: data = 8'hf9;
      17'd15687: data = 8'hdb;
      17'd15688: data = 8'h11;
      17'd15689: data = 8'h09;
      17'd15690: data = 8'hed;
      17'd15691: data = 8'h0c;
      17'd15692: data = 8'h0c;
      17'd15693: data = 8'hf1;
      17'd15694: data = 8'h0a;
      17'd15695: data = 8'hf6;
      17'd15696: data = 8'hf5;
      17'd15697: data = 8'h22;
      17'd15698: data = 8'hf6;
      17'd15699: data = 8'he5;
      17'd15700: data = 8'h11;
      17'd15701: data = 8'h04;
      17'd15702: data = 8'h00;
      17'd15703: data = 8'h13;
      17'd15704: data = 8'hf1;
      17'd15705: data = 8'he9;
      17'd15706: data = 8'h12;
      17'd15707: data = 8'h15;
      17'd15708: data = 8'hf4;
      17'd15709: data = 8'heb;
      17'd15710: data = 8'h05;
      17'd15711: data = 8'h0d;
      17'd15712: data = 8'hf6;
      17'd15713: data = 8'hf5;
      17'd15714: data = 8'hfe;
      17'd15715: data = 8'h01;
      17'd15716: data = 8'h00;
      17'd15717: data = 8'hfd;
      17'd15718: data = 8'h01;
      17'd15719: data = 8'hf1;
      17'd15720: data = 8'h01;
      17'd15721: data = 8'h0e;
      17'd15722: data = 8'hef;
      17'd15723: data = 8'hf1;
      17'd15724: data = 8'h0d;
      17'd15725: data = 8'hfa;
      17'd15726: data = 8'he7;
      17'd15727: data = 8'h01;
      17'd15728: data = 8'hf6;
      17'd15729: data = 8'h00;
      17'd15730: data = 8'h02;
      17'd15731: data = 8'heb;
      17'd15732: data = 8'h02;
      17'd15733: data = 8'h04;
      17'd15734: data = 8'he7;
      17'd15735: data = 8'hf6;
      17'd15736: data = 8'h13;
      17'd15737: data = 8'h04;
      17'd15738: data = 8'he5;
      17'd15739: data = 8'hfa;
      17'd15740: data = 8'h04;
      17'd15741: data = 8'hfc;
      17'd15742: data = 8'hfd;
      17'd15743: data = 8'hec;
      17'd15744: data = 8'h04;
      17'd15745: data = 8'h12;
      17'd15746: data = 8'hda;
      17'd15747: data = 8'hef;
      17'd15748: data = 8'h1e;
      17'd15749: data = 8'h04;
      17'd15750: data = 8'hf4;
      17'd15751: data = 8'hfc;
      17'd15752: data = 8'hfa;
      17'd15753: data = 8'h0d;
      17'd15754: data = 8'hf6;
      17'd15755: data = 8'heb;
      17'd15756: data = 8'h13;
      17'd15757: data = 8'h02;
      17'd15758: data = 8'hf2;
      17'd15759: data = 8'h00;
      17'd15760: data = 8'hf6;
      17'd15761: data = 8'h06;
      17'd15762: data = 8'h06;
      17'd15763: data = 8'he9;
      17'd15764: data = 8'h0c;
      17'd15765: data = 8'h06;
      17'd15766: data = 8'hf1;
      17'd15767: data = 8'h0e;
      17'd15768: data = 8'hfc;
      17'd15769: data = 8'he2;
      17'd15770: data = 8'h1a;
      17'd15771: data = 8'h0e;
      17'd15772: data = 8'hd6;
      17'd15773: data = 8'h09;
      17'd15774: data = 8'h15;
      17'd15775: data = 8'he7;
      17'd15776: data = 8'hf5;
      17'd15777: data = 8'h0e;
      17'd15778: data = 8'h05;
      17'd15779: data = 8'h06;
      17'd15780: data = 8'hf4;
      17'd15781: data = 8'he7;
      17'd15782: data = 8'hfe;
      17'd15783: data = 8'h11;
      17'd15784: data = 8'h09;
      17'd15785: data = 8'hf5;
      17'd15786: data = 8'hf1;
      17'd15787: data = 8'hf6;
      17'd15788: data = 8'hfe;
      17'd15789: data = 8'h0d;
      17'd15790: data = 8'hfd;
      17'd15791: data = 8'hfa;
      17'd15792: data = 8'h00;
      17'd15793: data = 8'hf6;
      17'd15794: data = 8'h04;
      17'd15795: data = 8'h04;
      17'd15796: data = 8'hf6;
      17'd15797: data = 8'h04;
      17'd15798: data = 8'hf9;
      17'd15799: data = 8'heb;
      17'd15800: data = 8'h0c;
      17'd15801: data = 8'h0c;
      17'd15802: data = 8'hed;
      17'd15803: data = 8'hf1;
      17'd15804: data = 8'h01;
      17'd15805: data = 8'h0c;
      17'd15806: data = 8'h00;
      17'd15807: data = 8'hf1;
      17'd15808: data = 8'hf5;
      17'd15809: data = 8'h05;
      17'd15810: data = 8'h0a;
      17'd15811: data = 8'hf2;
      17'd15812: data = 8'h04;
      17'd15813: data = 8'h06;
      17'd15814: data = 8'he3;
      17'd15815: data = 8'h01;
      17'd15816: data = 8'h1f;
      17'd15817: data = 8'he5;
      17'd15818: data = 8'hef;
      17'd15819: data = 8'h24;
      17'd15820: data = 8'he4;
      17'd15821: data = 8'he3;
      17'd15822: data = 8'h29;
      17'd15823: data = 8'h05;
      17'd15824: data = 8'he7;
      17'd15825: data = 8'h06;
      17'd15826: data = 8'hfd;
      17'd15827: data = 8'hf2;
      17'd15828: data = 8'h09;
      17'd15829: data = 8'h11;
      17'd15830: data = 8'h00;
      17'd15831: data = 8'hf2;
      17'd15832: data = 8'h01;
      17'd15833: data = 8'h0d;
      17'd15834: data = 8'hfa;
      17'd15835: data = 8'h05;
      17'd15836: data = 8'h13;
      17'd15837: data = 8'hef;
      17'd15838: data = 8'hfe;
      17'd15839: data = 8'h1a;
      17'd15840: data = 8'h05;
      17'd15841: data = 8'hfe;
      17'd15842: data = 8'h06;
      17'd15843: data = 8'h04;
      17'd15844: data = 8'hfc;
      17'd15845: data = 8'h0c;
      17'd15846: data = 8'h02;
      17'd15847: data = 8'hfe;
      17'd15848: data = 8'h15;
      17'd15849: data = 8'hfc;
      17'd15850: data = 8'hf5;
      17'd15851: data = 8'h1c;
      17'd15852: data = 8'h05;
      17'd15853: data = 8'hed;
      17'd15854: data = 8'h19;
      17'd15855: data = 8'h13;
      17'd15856: data = 8'hed;
      17'd15857: data = 8'h02;
      17'd15858: data = 8'h1b;
      17'd15859: data = 8'hf6;
      17'd15860: data = 8'hfc;
      17'd15861: data = 8'h13;
      17'd15862: data = 8'hfe;
      17'd15863: data = 8'hfa;
      17'd15864: data = 8'h0c;
      17'd15865: data = 8'h09;
      17'd15866: data = 8'hf9;
      17'd15867: data = 8'h01;
      17'd15868: data = 8'h11;
      17'd15869: data = 8'h02;
      17'd15870: data = 8'hf9;
      17'd15871: data = 8'h04;
      17'd15872: data = 8'h04;
      17'd15873: data = 8'hf2;
      17'd15874: data = 8'h09;
      17'd15875: data = 8'h13;
      17'd15876: data = 8'hec;
      17'd15877: data = 8'hed;
      17'd15878: data = 8'h12;
      17'd15879: data = 8'h04;
      17'd15880: data = 8'hec;
      17'd15881: data = 8'h05;
      17'd15882: data = 8'hfc;
      17'd15883: data = 8'hf9;
      17'd15884: data = 8'h16;
      17'd15885: data = 8'hf5;
      17'd15886: data = 8'hf4;
      17'd15887: data = 8'h0a;
      17'd15888: data = 8'hf6;
      17'd15889: data = 8'hf2;
      17'd15890: data = 8'h0c;
      17'd15891: data = 8'h00;
      17'd15892: data = 8'heb;
      17'd15893: data = 8'h04;
      17'd15894: data = 8'hf9;
      17'd15895: data = 8'hf6;
      17'd15896: data = 8'h12;
      17'd15897: data = 8'he9;
      17'd15898: data = 8'hf2;
      17'd15899: data = 8'h13;
      17'd15900: data = 8'heb;
      17'd15901: data = 8'hfc;
      17'd15902: data = 8'h13;
      17'd15903: data = 8'he9;
      17'd15904: data = 8'hfa;
      17'd15905: data = 8'h0c;
      17'd15906: data = 8'hf4;
      17'd15907: data = 8'h02;
      17'd15908: data = 8'h01;
      17'd15909: data = 8'hf2;
      17'd15910: data = 8'h09;
      17'd15911: data = 8'h06;
      17'd15912: data = 8'hf6;
      17'd15913: data = 8'h05;
      17'd15914: data = 8'h00;
      17'd15915: data = 8'heb;
      17'd15916: data = 8'h06;
      17'd15917: data = 8'h1e;
      17'd15918: data = 8'hec;
      17'd15919: data = 8'hf1;
      17'd15920: data = 8'h11;
      17'd15921: data = 8'hf6;
      17'd15922: data = 8'hf5;
      17'd15923: data = 8'h13;
      17'd15924: data = 8'h0c;
      17'd15925: data = 8'heb;
      17'd15926: data = 8'hfd;
      17'd15927: data = 8'h11;
      17'd15928: data = 8'h09;
      17'd15929: data = 8'hfe;
      17'd15930: data = 8'hfd;
      17'd15931: data = 8'h04;
      17'd15932: data = 8'h00;
      17'd15933: data = 8'hfd;
      17'd15934: data = 8'h06;
      17'd15935: data = 8'h0e;
      17'd15936: data = 8'hfe;
      17'd15937: data = 8'hf4;
      17'd15938: data = 8'h02;
      17'd15939: data = 8'h09;
      17'd15940: data = 8'hfc;
      17'd15941: data = 8'h05;
      17'd15942: data = 8'h06;
      17'd15943: data = 8'hfc;
      17'd15944: data = 8'hfd;
      17'd15945: data = 8'hfd;
      17'd15946: data = 8'h01;
      17'd15947: data = 8'h09;
      17'd15948: data = 8'h04;
      17'd15949: data = 8'hf5;
      17'd15950: data = 8'heb;
      17'd15951: data = 8'h01;
      17'd15952: data = 8'h11;
      17'd15953: data = 8'hfa;
      17'd15954: data = 8'hf2;
      17'd15955: data = 8'hfe;
      17'd15956: data = 8'h09;
      17'd15957: data = 8'hfa;
      17'd15958: data = 8'hf4;
      17'd15959: data = 8'h00;
      17'd15960: data = 8'h02;
      17'd15961: data = 8'hf9;
      17'd15962: data = 8'he9;
      17'd15963: data = 8'h02;
      17'd15964: data = 8'h06;
      17'd15965: data = 8'he4;
      17'd15966: data = 8'hfa;
      17'd15967: data = 8'h19;
      17'd15968: data = 8'hf1;
      17'd15969: data = 8'he4;
      17'd15970: data = 8'h09;
      17'd15971: data = 8'h05;
      17'd15972: data = 8'hf6;
      17'd15973: data = 8'h09;
      17'd15974: data = 8'hfd;
      17'd15975: data = 8'he5;
      17'd15976: data = 8'hfc;
      17'd15977: data = 8'h13;
      17'd15978: data = 8'h02;
      17'd15979: data = 8'hf5;
      17'd15980: data = 8'hf6;
      17'd15981: data = 8'hfc;
      17'd15982: data = 8'h06;
      17'd15983: data = 8'h0a;
      17'd15984: data = 8'h01;
      17'd15985: data = 8'hfa;
      17'd15986: data = 8'hfc;
      17'd15987: data = 8'h09;
      17'd15988: data = 8'h0e;
      17'd15989: data = 8'hf5;
      17'd15990: data = 8'hf5;
      17'd15991: data = 8'h06;
      17'd15992: data = 8'h04;
      17'd15993: data = 8'h0e;
      17'd15994: data = 8'hfd;
      17'd15995: data = 8'hf4;
      17'd15996: data = 8'h01;
      17'd15997: data = 8'h04;
      17'd15998: data = 8'h19;
      17'd15999: data = 8'h0a;
      17'd16000: data = 8'he9;
      17'd16001: data = 8'hfd;
      17'd16002: data = 8'h0e;
      17'd16003: data = 8'hf9;
      17'd16004: data = 8'h02;
      17'd16005: data = 8'h13;
      17'd16006: data = 8'hf4;
      17'd16007: data = 8'hf1;
      17'd16008: data = 8'h0c;
      17'd16009: data = 8'h0d;
      17'd16010: data = 8'hfc;
      17'd16011: data = 8'hf2;
      17'd16012: data = 8'h0c;
      17'd16013: data = 8'h06;
      17'd16014: data = 8'hf4;
      17'd16015: data = 8'h0d;
      17'd16016: data = 8'hfe;
      17'd16017: data = 8'hef;
      17'd16018: data = 8'h0a;
      17'd16019: data = 8'h04;
      17'd16020: data = 8'hf4;
      17'd16021: data = 8'hfd;
      17'd16022: data = 8'h02;
      17'd16023: data = 8'hf6;
      17'd16024: data = 8'h00;
      17'd16025: data = 8'hfe;
      17'd16026: data = 8'hfa;
      17'd16027: data = 8'h09;
      17'd16028: data = 8'hf2;
      17'd16029: data = 8'hf4;
      17'd16030: data = 8'h0a;
      17'd16031: data = 8'hf4;
      17'd16032: data = 8'hed;
      17'd16033: data = 8'h0d;
      17'd16034: data = 8'hfe;
      17'd16035: data = 8'he9;
      17'd16036: data = 8'h0c;
      17'd16037: data = 8'hf6;
      17'd16038: data = 8'heb;
      17'd16039: data = 8'h0d;
      17'd16040: data = 8'hfd;
      17'd16041: data = 8'hed;
      17'd16042: data = 8'h00;
      17'd16043: data = 8'h05;
      17'd16044: data = 8'hfa;
      17'd16045: data = 8'hec;
      17'd16046: data = 8'h00;
      17'd16047: data = 8'h0e;
      17'd16048: data = 8'hf9;
      17'd16049: data = 8'heb;
      17'd16050: data = 8'h05;
      17'd16051: data = 8'h0c;
      17'd16052: data = 8'hec;
      17'd16053: data = 8'hfc;
      17'd16054: data = 8'h0a;
      17'd16055: data = 8'hfd;
      17'd16056: data = 8'hfa;
      17'd16057: data = 8'h04;
      17'd16058: data = 8'h0a;
      17'd16059: data = 8'hfa;
      17'd16060: data = 8'h04;
      17'd16061: data = 8'h11;
      17'd16062: data = 8'hf6;
      17'd16063: data = 8'hf5;
      17'd16064: data = 8'h13;
      17'd16065: data = 8'h0d;
      17'd16066: data = 8'hed;
      17'd16067: data = 8'h06;
      17'd16068: data = 8'h19;
      17'd16069: data = 8'hf6;
      17'd16070: data = 8'hfc;
      17'd16071: data = 8'h15;
      17'd16072: data = 8'h11;
      17'd16073: data = 8'hfc;
      17'd16074: data = 8'hf9;
      17'd16075: data = 8'h11;
      17'd16076: data = 8'h05;
      17'd16077: data = 8'h04;
      17'd16078: data = 8'h11;
      17'd16079: data = 8'hfe;
      17'd16080: data = 8'hf9;
      17'd16081: data = 8'h04;
      17'd16082: data = 8'h0a;
      17'd16083: data = 8'h01;
      17'd16084: data = 8'h02;
      17'd16085: data = 8'h09;
      17'd16086: data = 8'h00;
      17'd16087: data = 8'hfa;
      17'd16088: data = 8'h02;
      17'd16089: data = 8'h12;
      17'd16090: data = 8'hfc;
      17'd16091: data = 8'hf6;
      17'd16092: data = 8'h11;
      17'd16093: data = 8'h05;
      17'd16094: data = 8'hf5;
      17'd16095: data = 8'h01;
      17'd16096: data = 8'h0e;
      17'd16097: data = 8'h00;
      17'd16098: data = 8'hed;
      17'd16099: data = 8'h01;
      17'd16100: data = 8'h05;
      17'd16101: data = 8'hfa;
      17'd16102: data = 8'hfe;
      17'd16103: data = 8'h04;
      17'd16104: data = 8'hf5;
      17'd16105: data = 8'hfe;
      17'd16106: data = 8'h0e;
      17'd16107: data = 8'hfc;
      17'd16108: data = 8'he9;
      17'd16109: data = 8'h06;
      17'd16110: data = 8'h0c;
      17'd16111: data = 8'hed;
      17'd16112: data = 8'hf4;
      17'd16113: data = 8'hfe;
      17'd16114: data = 8'hfa;
      17'd16115: data = 8'h00;
      17'd16116: data = 8'h01;
      17'd16117: data = 8'hf2;
      17'd16118: data = 8'hf5;
      17'd16119: data = 8'h05;
      17'd16120: data = 8'hfe;
      17'd16121: data = 8'hf9;
      17'd16122: data = 8'h01;
      17'd16123: data = 8'hfe;
      17'd16124: data = 8'hfa;
      17'd16125: data = 8'hf5;
      17'd16126: data = 8'hfa;
      17'd16127: data = 8'h02;
      17'd16128: data = 8'hf9;
      17'd16129: data = 8'hfa;
      17'd16130: data = 8'h00;
      17'd16131: data = 8'hf6;
      17'd16132: data = 8'hfc;
      17'd16133: data = 8'h02;
      17'd16134: data = 8'h01;
      17'd16135: data = 8'hfa;
      17'd16136: data = 8'hf4;
      17'd16137: data = 8'h01;
      17'd16138: data = 8'h05;
      17'd16139: data = 8'hfe;
      17'd16140: data = 8'hfe;
      17'd16141: data = 8'h02;
      17'd16142: data = 8'hf6;
      17'd16143: data = 8'hf6;
      17'd16144: data = 8'h11;
      17'd16145: data = 8'h01;
      17'd16146: data = 8'hfa;
      17'd16147: data = 8'h06;
      17'd16148: data = 8'hfa;
      17'd16149: data = 8'h05;
      17'd16150: data = 8'h13;
      17'd16151: data = 8'hfa;
      17'd16152: data = 8'hf6;
      17'd16153: data = 8'h0a;
      17'd16154: data = 8'h04;
      17'd16155: data = 8'h0c;
      17'd16156: data = 8'h04;
      17'd16157: data = 8'hf2;
      17'd16158: data = 8'h05;
      17'd16159: data = 8'h11;
      17'd16160: data = 8'h01;
      17'd16161: data = 8'hfd;
      17'd16162: data = 8'hf6;
      17'd16163: data = 8'hfd;
      17'd16164: data = 8'h0c;
      17'd16165: data = 8'h0a;
      17'd16166: data = 8'hfa;
      17'd16167: data = 8'hf5;
      17'd16168: data = 8'h05;
      17'd16169: data = 8'h02;
      17'd16170: data = 8'hf1;
      17'd16171: data = 8'h01;
      17'd16172: data = 8'h02;
      17'd16173: data = 8'hec;
      17'd16174: data = 8'h02;
      17'd16175: data = 8'h0e;
      17'd16176: data = 8'hec;
      17'd16177: data = 8'hed;
      17'd16178: data = 8'h09;
      17'd16179: data = 8'h05;
      17'd16180: data = 8'hf1;
      17'd16181: data = 8'hfe;
      17'd16182: data = 8'hf9;
      17'd16183: data = 8'he7;
      17'd16184: data = 8'h0c;
      17'd16185: data = 8'h0a;
      17'd16186: data = 8'he9;
      17'd16187: data = 8'hf6;
      17'd16188: data = 8'h09;
      17'd16189: data = 8'hfd;
      17'd16190: data = 8'hf5;
      17'd16191: data = 8'h00;
      17'd16192: data = 8'hfe;
      17'd16193: data = 8'hf9;
      17'd16194: data = 8'h02;
      17'd16195: data = 8'h05;
      17'd16196: data = 8'hf5;
      17'd16197: data = 8'h00;
      17'd16198: data = 8'h01;
      17'd16199: data = 8'hf5;
      17'd16200: data = 8'h05;
      17'd16201: data = 8'h04;
      17'd16202: data = 8'hf5;
      17'd16203: data = 8'h04;
      17'd16204: data = 8'h09;
      17'd16205: data = 8'h00;
      17'd16206: data = 8'h05;
      17'd16207: data = 8'h02;
      17'd16208: data = 8'hfc;
      17'd16209: data = 8'h02;
      17'd16210: data = 8'h09;
      17'd16211: data = 8'hfd;
      17'd16212: data = 8'hf5;
      17'd16213: data = 8'h05;
      17'd16214: data = 8'h11;
      17'd16215: data = 8'h06;
      17'd16216: data = 8'hfe;
      17'd16217: data = 8'hfc;
      17'd16218: data = 8'h06;
      17'd16219: data = 8'hfd;
      17'd16220: data = 8'hfc;
      17'd16221: data = 8'h16;
      17'd16222: data = 8'h02;
      17'd16223: data = 8'hef;
      17'd16224: data = 8'hfd;
      17'd16225: data = 8'h00;
      17'd16226: data = 8'h06;
      17'd16227: data = 8'h04;
      17'd16228: data = 8'hf6;
      17'd16229: data = 8'h00;
      17'd16230: data = 8'h06;
      17'd16231: data = 8'hf5;
      17'd16232: data = 8'hf6;
      17'd16233: data = 8'h09;
      17'd16234: data = 8'h06;
      17'd16235: data = 8'hfc;
      17'd16236: data = 8'hfa;
      17'd16237: data = 8'hfa;
      17'd16238: data = 8'h01;
      17'd16239: data = 8'h05;
      17'd16240: data = 8'hfd;
      17'd16241: data = 8'hfd;
      17'd16242: data = 8'hfe;
      17'd16243: data = 8'hf5;
      17'd16244: data = 8'hfe;
      17'd16245: data = 8'h01;
      17'd16246: data = 8'hf6;
      17'd16247: data = 8'hfe;
      17'd16248: data = 8'h00;
      17'd16249: data = 8'hfa;
      17'd16250: data = 8'hfc;
      17'd16251: data = 8'hf6;
      17'd16252: data = 8'hf6;
      17'd16253: data = 8'hfe;
      17'd16254: data = 8'h02;
      17'd16255: data = 8'hfd;
      17'd16256: data = 8'hf9;
      17'd16257: data = 8'hf2;
      17'd16258: data = 8'hf6;
      17'd16259: data = 8'h02;
      17'd16260: data = 8'h05;
      17'd16261: data = 8'h00;
      17'd16262: data = 8'hf2;
      17'd16263: data = 8'hf9;
      17'd16264: data = 8'h00;
      17'd16265: data = 8'hfc;
      17'd16266: data = 8'hfe;
      17'd16267: data = 8'h09;
      17'd16268: data = 8'h01;
      17'd16269: data = 8'hf1;
      17'd16270: data = 8'hf2;
      17'd16271: data = 8'h00;
      17'd16272: data = 8'h02;
      17'd16273: data = 8'hfe;
      17'd16274: data = 8'h04;
      17'd16275: data = 8'hfe;
      17'd16276: data = 8'hf1;
      17'd16277: data = 8'hfe;
      17'd16278: data = 8'h0a;
      17'd16279: data = 8'h04;
      17'd16280: data = 8'hfd;
      17'd16281: data = 8'hfd;
      17'd16282: data = 8'hfc;
      17'd16283: data = 8'hfd;
      17'd16284: data = 8'h0a;
      17'd16285: data = 8'h05;
      17'd16286: data = 8'h00;
      17'd16287: data = 8'h01;
      17'd16288: data = 8'hfe;
      17'd16289: data = 8'h09;
      17'd16290: data = 8'h09;
      17'd16291: data = 8'hfd;
      17'd16292: data = 8'hfe;
      17'd16293: data = 8'h0a;
      17'd16294: data = 8'h0d;
      17'd16295: data = 8'h02;
      17'd16296: data = 8'hfc;
      17'd16297: data = 8'h01;
      17'd16298: data = 8'h06;
      17'd16299: data = 8'h05;
      17'd16300: data = 8'h04;
      17'd16301: data = 8'h04;
      17'd16302: data = 8'h00;
      17'd16303: data = 8'hfd;
      17'd16304: data = 8'h05;
      17'd16305: data = 8'h0a;
      17'd16306: data = 8'h02;
      17'd16307: data = 8'hfd;
      17'd16308: data = 8'h01;
      17'd16309: data = 8'h02;
      17'd16310: data = 8'h02;
      17'd16311: data = 8'h01;
      17'd16312: data = 8'h01;
      17'd16313: data = 8'h09;
      17'd16314: data = 8'h09;
      17'd16315: data = 8'hfa;
      17'd16316: data = 8'hfd;
      17'd16317: data = 8'h0d;
      17'd16318: data = 8'h04;
      17'd16319: data = 8'hfa;
      17'd16320: data = 8'h04;
      17'd16321: data = 8'h04;
      17'd16322: data = 8'hfc;
      17'd16323: data = 8'h04;
      17'd16324: data = 8'h04;
      17'd16325: data = 8'h00;
      17'd16326: data = 8'hfd;
      17'd16327: data = 8'h01;
      17'd16328: data = 8'h00;
      17'd16329: data = 8'hfe;
      17'd16330: data = 8'h02;
      17'd16331: data = 8'h00;
      17'd16332: data = 8'h01;
      17'd16333: data = 8'h01;
      17'd16334: data = 8'h01;
      17'd16335: data = 8'hfa;
      17'd16336: data = 8'hfa;
      17'd16337: data = 8'h01;
      17'd16338: data = 8'h02;
      17'd16339: data = 8'hfd;
      17'd16340: data = 8'hfe;
      17'd16341: data = 8'hfe;
      17'd16342: data = 8'h00;
      17'd16343: data = 8'h05;
      17'd16344: data = 8'h00;
      17'd16345: data = 8'hf5;
      17'd16346: data = 8'hfd;
      17'd16347: data = 8'h00;
      17'd16348: data = 8'h00;
      17'd16349: data = 8'h00;
      17'd16350: data = 8'hfa;
      17'd16351: data = 8'hf9;
      17'd16352: data = 8'hfe;
      17'd16353: data = 8'hfe;
      17'd16354: data = 8'hf9;
      17'd16355: data = 8'hfe;
      17'd16356: data = 8'h02;
      17'd16357: data = 8'hfa;
      17'd16358: data = 8'hf4;
      17'd16359: data = 8'h05;
      17'd16360: data = 8'h06;
      17'd16361: data = 8'hf6;
      17'd16362: data = 8'hfa;
      17'd16363: data = 8'hf9;
      17'd16364: data = 8'hf9;
      17'd16365: data = 8'hfa;
      17'd16366: data = 8'hfe;
      17'd16367: data = 8'h02;
      17'd16368: data = 8'hfe;
      17'd16369: data = 8'hfd;
      17'd16370: data = 8'hf6;
      17'd16371: data = 8'hfe;
      17'd16372: data = 8'h09;
      17'd16373: data = 8'hfd;
      17'd16374: data = 8'hf6;
      17'd16375: data = 8'h02;
      17'd16376: data = 8'h04;
      17'd16377: data = 8'hfe;
      17'd16378: data = 8'h04;
      17'd16379: data = 8'hf5;
      17'd16380: data = 8'hf2;
      17'd16381: data = 8'h0e;
      17'd16382: data = 8'h09;
      17'd16383: data = 8'hf2;
      17'd16384: data = 8'hfa;
      17'd16385: data = 8'h05;
      17'd16386: data = 8'h05;
      17'd16387: data = 8'h05;
      17'd16388: data = 8'h01;
      17'd16389: data = 8'hfd;
      17'd16390: data = 8'hfe;
      17'd16391: data = 8'hfc;
      17'd16392: data = 8'hfc;
      17'd16393: data = 8'h04;
      17'd16394: data = 8'h05;
      17'd16395: data = 8'hfc;
      17'd16396: data = 8'hfc;
      17'd16397: data = 8'h01;
      17'd16398: data = 8'h00;
      17'd16399: data = 8'hf9;
      17'd16400: data = 8'hfd;
      17'd16401: data = 8'h04;
      17'd16402: data = 8'h00;
      17'd16403: data = 8'hfc;
      17'd16404: data = 8'hfe;
      17'd16405: data = 8'hfc;
      17'd16406: data = 8'hfc;
      17'd16407: data = 8'h01;
      17'd16408: data = 8'hf9;
      17'd16409: data = 8'hf4;
      17'd16410: data = 8'hfd;
      17'd16411: data = 8'h01;
      17'd16412: data = 8'hfd;
      17'd16413: data = 8'hfa;
      17'd16414: data = 8'h00;
      17'd16415: data = 8'h01;
      17'd16416: data = 8'hfd;
      17'd16417: data = 8'hfc;
      17'd16418: data = 8'hf9;
      17'd16419: data = 8'hf9;
      17'd16420: data = 8'hfc;
      17'd16421: data = 8'h00;
      17'd16422: data = 8'hfe;
      17'd16423: data = 8'hf5;
      17'd16424: data = 8'hfc;
      17'd16425: data = 8'h02;
      17'd16426: data = 8'hfa;
      17'd16427: data = 8'h00;
      17'd16428: data = 8'h04;
      17'd16429: data = 8'hf6;
      17'd16430: data = 8'hfc;
      17'd16431: data = 8'h01;
      17'd16432: data = 8'hfe;
      17'd16433: data = 8'h00;
      17'd16434: data = 8'h01;
      17'd16435: data = 8'hfd;
      17'd16436: data = 8'hfd;
      17'd16437: data = 8'hfc;
      17'd16438: data = 8'hfe;
      17'd16439: data = 8'h06;
      17'd16440: data = 8'h02;
      17'd16441: data = 8'h05;
      17'd16442: data = 8'h04;
      17'd16443: data = 8'hfc;
      17'd16444: data = 8'hfe;
      17'd16445: data = 8'h02;
      17'd16446: data = 8'h04;
      17'd16447: data = 8'h04;
      17'd16448: data = 8'h02;
      17'd16449: data = 8'hf9;
      17'd16450: data = 8'hfe;
      17'd16451: data = 8'h04;
      17'd16452: data = 8'hfd;
      17'd16453: data = 8'h00;
      17'd16454: data = 8'h05;
      17'd16455: data = 8'hfe;
      17'd16456: data = 8'h01;
      17'd16457: data = 8'h04;
      17'd16458: data = 8'hfe;
      17'd16459: data = 8'h02;
      17'd16460: data = 8'h04;
      17'd16461: data = 8'hfd;
      17'd16462: data = 8'hfe;
      17'd16463: data = 8'hfe;
      17'd16464: data = 8'hfa;
      17'd16465: data = 8'h04;
      17'd16466: data = 8'h04;
      17'd16467: data = 8'hfd;
      17'd16468: data = 8'h00;
      17'd16469: data = 8'hfd;
      17'd16470: data = 8'hfc;
      17'd16471: data = 8'h02;
      17'd16472: data = 8'hfe;
      17'd16473: data = 8'hfc;
      17'd16474: data = 8'h00;
      17'd16475: data = 8'hfd;
      17'd16476: data = 8'hf9;
      17'd16477: data = 8'hfd;
      17'd16478: data = 8'hf9;
      17'd16479: data = 8'hf5;
      17'd16480: data = 8'hfe;
      17'd16481: data = 8'hfc;
      17'd16482: data = 8'hf5;
      17'd16483: data = 8'hfc;
      17'd16484: data = 8'hfe;
      17'd16485: data = 8'hfa;
      17'd16486: data = 8'hf6;
      17'd16487: data = 8'hfa;
      17'd16488: data = 8'hfc;
      17'd16489: data = 8'hf2;
      17'd16490: data = 8'hf1;
      17'd16491: data = 8'hfd;
      17'd16492: data = 8'hfc;
      17'd16493: data = 8'hf4;
      17'd16494: data = 8'hfe;
      17'd16495: data = 8'hfe;
      17'd16496: data = 8'hf4;
      17'd16497: data = 8'hfd;
      17'd16498: data = 8'h00;
      17'd16499: data = 8'hfc;
      17'd16500: data = 8'hfe;
      17'd16501: data = 8'h00;
      17'd16502: data = 8'hfd;
      17'd16503: data = 8'h00;
      17'd16504: data = 8'h02;
      17'd16505: data = 8'h01;
      17'd16506: data = 8'h00;
      17'd16507: data = 8'h02;
      17'd16508: data = 8'h02;
      17'd16509: data = 8'h04;
      17'd16510: data = 8'h05;
      17'd16511: data = 8'h04;
      17'd16512: data = 8'h0a;
      17'd16513: data = 8'h06;
      17'd16514: data = 8'h00;
      17'd16515: data = 8'h06;
      17'd16516: data = 8'h0a;
      17'd16517: data = 8'h01;
      17'd16518: data = 8'h04;
      17'd16519: data = 8'h06;
      17'd16520: data = 8'h04;
      17'd16521: data = 8'h04;
      17'd16522: data = 8'h09;
      17'd16523: data = 8'h09;
      17'd16524: data = 8'h04;
      17'd16525: data = 8'h05;
      17'd16526: data = 8'h0a;
      17'd16527: data = 8'h0a;
      17'd16528: data = 8'h05;
      17'd16529: data = 8'h04;
      17'd16530: data = 8'h04;
      17'd16531: data = 8'h02;
      17'd16532: data = 8'h01;
      17'd16533: data = 8'h00;
      17'd16534: data = 8'h02;
      17'd16535: data = 8'h00;
      17'd16536: data = 8'hfd;
      17'd16537: data = 8'h00;
      17'd16538: data = 8'h00;
      17'd16539: data = 8'hfc;
      17'd16540: data = 8'hf9;
      17'd16541: data = 8'hfc;
      17'd16542: data = 8'hfe;
      17'd16543: data = 8'h02;
      17'd16544: data = 8'hfd;
      17'd16545: data = 8'hf6;
      17'd16546: data = 8'hfc;
      17'd16547: data = 8'hfe;
      17'd16548: data = 8'hfd;
      17'd16549: data = 8'hfe;
      17'd16550: data = 8'hfa;
      17'd16551: data = 8'hf6;
      17'd16552: data = 8'hfe;
      17'd16553: data = 8'h01;
      17'd16554: data = 8'hfe;
      17'd16555: data = 8'h00;
      17'd16556: data = 8'h01;
      17'd16557: data = 8'hfe;
      17'd16558: data = 8'hfe;
      17'd16559: data = 8'h00;
      17'd16560: data = 8'h02;
      17'd16561: data = 8'h04;
      17'd16562: data = 8'h02;
      17'd16563: data = 8'h02;
      17'd16564: data = 8'h05;
      17'd16565: data = 8'h02;
      17'd16566: data = 8'h02;
      17'd16567: data = 8'h06;
      17'd16568: data = 8'h09;
      17'd16569: data = 8'h06;
      17'd16570: data = 8'h06;
      17'd16571: data = 8'h05;
      17'd16572: data = 8'h06;
      17'd16573: data = 8'h0c;
      17'd16574: data = 8'h06;
      17'd16575: data = 8'h04;
      17'd16576: data = 8'h06;
      17'd16577: data = 8'h05;
      17'd16578: data = 8'h02;
      17'd16579: data = 8'h05;
      17'd16580: data = 8'h04;
      17'd16581: data = 8'h01;
      17'd16582: data = 8'h02;
      17'd16583: data = 8'h02;
      17'd16584: data = 8'h04;
      17'd16585: data = 8'h05;
      17'd16586: data = 8'h00;
      17'd16587: data = 8'hfd;
      17'd16588: data = 8'h01;
      17'd16589: data = 8'h04;
      17'd16590: data = 8'h02;
      17'd16591: data = 8'h00;
      17'd16592: data = 8'h00;
      17'd16593: data = 8'h00;
      17'd16594: data = 8'h00;
      17'd16595: data = 8'hfc;
      17'd16596: data = 8'hfd;
      17'd16597: data = 8'h00;
      17'd16598: data = 8'hfd;
      17'd16599: data = 8'hfc;
      17'd16600: data = 8'hfe;
      17'd16601: data = 8'hfe;
      17'd16602: data = 8'hf6;
      17'd16603: data = 8'hf4;
      17'd16604: data = 8'h01;
      17'd16605: data = 8'h04;
      17'd16606: data = 8'hfd;
      17'd16607: data = 8'hf9;
      17'd16608: data = 8'hf9;
      17'd16609: data = 8'hfe;
      17'd16610: data = 8'hfe;
      17'd16611: data = 8'hfa;
      17'd16612: data = 8'hfa;
      17'd16613: data = 8'h01;
      17'd16614: data = 8'hfe;
      17'd16615: data = 8'hf6;
      17'd16616: data = 8'hfd;
      17'd16617: data = 8'hfa;
      17'd16618: data = 8'hf6;
      17'd16619: data = 8'h02;
      17'd16620: data = 8'hfc;
      17'd16621: data = 8'hf1;
      17'd16622: data = 8'hfc;
      17'd16623: data = 8'h02;
      17'd16624: data = 8'hf5;
      17'd16625: data = 8'hfd;
      17'd16626: data = 8'h06;
      17'd16627: data = 8'hfa;
      17'd16628: data = 8'hf2;
      17'd16629: data = 8'hf4;
      17'd16630: data = 8'h00;
      17'd16631: data = 8'hfc;
      17'd16632: data = 8'hf5;
      17'd16633: data = 8'hf4;
      17'd16634: data = 8'hfa;
      17'd16635: data = 8'hfc;
      17'd16636: data = 8'hf1;
      17'd16637: data = 8'hf4;
      17'd16638: data = 8'hfc;
      17'd16639: data = 8'hfc;
      17'd16640: data = 8'hf5;
      17'd16641: data = 8'hfa;
      17'd16642: data = 8'hf6;
      17'd16643: data = 8'hed;
      17'd16644: data = 8'hf9;
      17'd16645: data = 8'hfa;
      17'd16646: data = 8'hf5;
      17'd16647: data = 8'hf6;
      17'd16648: data = 8'hfa;
      17'd16649: data = 8'hfc;
      17'd16650: data = 8'hf1;
      17'd16651: data = 8'hfc;
      17'd16652: data = 8'hfc;
      17'd16653: data = 8'hef;
      17'd16654: data = 8'hf5;
      17'd16655: data = 8'hf6;
      17'd16656: data = 8'hfa;
      17'd16657: data = 8'hfe;
      17'd16658: data = 8'h04;
      17'd16659: data = 8'hef;
      17'd16660: data = 8'hed;
      17'd16661: data = 8'hfc;
      17'd16662: data = 8'hef;
      17'd16663: data = 8'hf1;
      17'd16664: data = 8'h00;
      17'd16665: data = 8'h06;
      17'd16666: data = 8'h05;
      17'd16667: data = 8'h0d;
      17'd16668: data = 8'h09;
      17'd16669: data = 8'h01;
      17'd16670: data = 8'h0c;
      17'd16671: data = 8'h06;
      17'd16672: data = 8'hfc;
      17'd16673: data = 8'h0e;
      17'd16674: data = 8'h16;
      17'd16675: data = 8'h02;
      17'd16676: data = 8'h09;
      17'd16677: data = 8'h11;
      17'd16678: data = 8'h04;
      17'd16679: data = 8'h0c;
      17'd16680: data = 8'h19;
      17'd16681: data = 8'h0a;
      17'd16682: data = 8'h09;
      17'd16683: data = 8'h12;
      17'd16684: data = 8'h11;
      17'd16685: data = 8'h0c;
      17'd16686: data = 8'h15;
      17'd16687: data = 8'h15;
      17'd16688: data = 8'h04;
      17'd16689: data = 8'hfe;
      17'd16690: data = 8'hfe;
      17'd16691: data = 8'hfe;
      17'd16692: data = 8'h02;
      17'd16693: data = 8'h00;
      17'd16694: data = 8'h00;
      17'd16695: data = 8'h0a;
      17'd16696: data = 8'h02;
      17'd16697: data = 8'hfa;
      17'd16698: data = 8'hfd;
      17'd16699: data = 8'hfd;
      17'd16700: data = 8'hfc;
      17'd16701: data = 8'hfc;
      17'd16702: data = 8'hf9;
      17'd16703: data = 8'hf6;
      17'd16704: data = 8'hfa;
      17'd16705: data = 8'hf4;
      17'd16706: data = 8'hec;
      17'd16707: data = 8'hf4;
      17'd16708: data = 8'hf4;
      17'd16709: data = 8'heb;
      17'd16710: data = 8'hec;
      17'd16711: data = 8'hef;
      17'd16712: data = 8'hed;
      17'd16713: data = 8'hf2;
      17'd16714: data = 8'hf1;
      17'd16715: data = 8'hf1;
      17'd16716: data = 8'hf1;
      17'd16717: data = 8'hec;
      17'd16718: data = 8'he9;
      17'd16719: data = 8'he7;
      17'd16720: data = 8'he9;
      17'd16721: data = 8'hef;
      17'd16722: data = 8'hf6;
      17'd16723: data = 8'hf5;
      17'd16724: data = 8'hf6;
      17'd16725: data = 8'hfa;
      17'd16726: data = 8'hfe;
      17'd16727: data = 8'h00;
      17'd16728: data = 8'h04;
      17'd16729: data = 8'h0e;
      17'd16730: data = 8'h0e;
      17'd16731: data = 8'h0e;
      17'd16732: data = 8'h11;
      17'd16733: data = 8'h16;
      17'd16734: data = 8'h1a;
      17'd16735: data = 8'h1a;
      17'd16736: data = 8'h1c;
      17'd16737: data = 8'h1e;
      17'd16738: data = 8'h24;
      17'd16739: data = 8'h27;
      17'd16740: data = 8'h27;
      17'd16741: data = 8'h2b;
      17'd16742: data = 8'h31;
      17'd16743: data = 8'h31;
      17'd16744: data = 8'h2b;
      17'd16745: data = 8'h2c;
      17'd16746: data = 8'h2c;
      17'd16747: data = 8'h22;
      17'd16748: data = 8'h1b;
      17'd16749: data = 8'h22;
      17'd16750: data = 8'h1c;
      17'd16751: data = 8'h19;
      17'd16752: data = 8'h16;
      17'd16753: data = 8'h13;
      17'd16754: data = 8'h16;
      17'd16755: data = 8'h13;
      17'd16756: data = 8'h13;
      17'd16757: data = 8'h11;
      17'd16758: data = 8'h0d;
      17'd16759: data = 8'h0a;
      17'd16760: data = 8'h0a;
      17'd16761: data = 8'h06;
      17'd16762: data = 8'hfd;
      17'd16763: data = 8'hfc;
      17'd16764: data = 8'hf9;
      17'd16765: data = 8'hf5;
      17'd16766: data = 8'hf2;
      17'd16767: data = 8'hed;
      17'd16768: data = 8'hef;
      17'd16769: data = 8'hef;
      17'd16770: data = 8'hec;
      17'd16771: data = 8'hed;
      17'd16772: data = 8'hef;
      17'd16773: data = 8'he9;
      17'd16774: data = 8'he7;
      17'd16775: data = 8'he7;
      17'd16776: data = 8'he3;
      17'd16777: data = 8'he2;
      17'd16778: data = 8'he3;
      17'd16779: data = 8'he3;
      17'd16780: data = 8'he2;
      17'd16781: data = 8'he0;
      17'd16782: data = 8'he0;
      17'd16783: data = 8'he5;
      17'd16784: data = 8'heb;
      17'd16785: data = 8'he9;
      17'd16786: data = 8'hec;
      17'd16787: data = 8'hed;
      17'd16788: data = 8'hec;
      17'd16789: data = 8'hed;
      17'd16790: data = 8'hef;
      17'd16791: data = 8'hf1;
      17'd16792: data = 8'hf2;
      17'd16793: data = 8'hed;
      17'd16794: data = 8'heb;
      17'd16795: data = 8'hed;
      17'd16796: data = 8'hf4;
      17'd16797: data = 8'hf6;
      17'd16798: data = 8'hf4;
      17'd16799: data = 8'hf2;
      17'd16800: data = 8'hf4;
      17'd16801: data = 8'hf6;
      17'd16802: data = 8'hf9;
      17'd16803: data = 8'hf5;
      17'd16804: data = 8'hf1;
      17'd16805: data = 8'hf2;
      17'd16806: data = 8'hf6;
      17'd16807: data = 8'hf5;
      17'd16808: data = 8'hf2;
      17'd16809: data = 8'hf4;
      17'd16810: data = 8'hf1;
      17'd16811: data = 8'hf1;
      17'd16812: data = 8'hf4;
      17'd16813: data = 8'hf6;
      17'd16814: data = 8'hf4;
      17'd16815: data = 8'hf4;
      17'd16816: data = 8'hfa;
      17'd16817: data = 8'hfa;
      17'd16818: data = 8'hf6;
      17'd16819: data = 8'hf4;
      17'd16820: data = 8'hf9;
      17'd16821: data = 8'hf6;
      17'd16822: data = 8'hf1;
      17'd16823: data = 8'hf9;
      17'd16824: data = 8'hfc;
      17'd16825: data = 8'hf4;
      17'd16826: data = 8'hf2;
      17'd16827: data = 8'hfa;
      17'd16828: data = 8'hfc;
      17'd16829: data = 8'hf5;
      17'd16830: data = 8'hfd;
      17'd16831: data = 8'hfe;
      17'd16832: data = 8'hfa;
      17'd16833: data = 8'hfe;
      17'd16834: data = 8'h02;
      17'd16835: data = 8'h04;
      17'd16836: data = 8'hfa;
      17'd16837: data = 8'hfc;
      17'd16838: data = 8'h01;
      17'd16839: data = 8'h01;
      17'd16840: data = 8'h02;
      17'd16841: data = 8'h04;
      17'd16842: data = 8'h0e;
      17'd16843: data = 8'h0c;
      17'd16844: data = 8'h04;
      17'd16845: data = 8'h05;
      17'd16846: data = 8'h06;
      17'd16847: data = 8'h0e;
      17'd16848: data = 8'h09;
      17'd16849: data = 8'hfe;
      17'd16850: data = 8'h09;
      17'd16851: data = 8'h0a;
      17'd16852: data = 8'h09;
      17'd16853: data = 8'h02;
      17'd16854: data = 8'h09;
      17'd16855: data = 8'h0e;
      17'd16856: data = 8'hfa;
      17'd16857: data = 8'h04;
      17'd16858: data = 8'h0c;
      17'd16859: data = 8'h04;
      17'd16860: data = 8'h12;
      17'd16861: data = 8'h0e;
      17'd16862: data = 8'hfd;
      17'd16863: data = 8'hfa;
      17'd16864: data = 8'hfd;
      17'd16865: data = 8'hf5;
      17'd16866: data = 8'hfa;
      17'd16867: data = 8'h0e;
      17'd16868: data = 8'h04;
      17'd16869: data = 8'hf2;
      17'd16870: data = 8'h00;
      17'd16871: data = 8'h02;
      17'd16872: data = 8'he5;
      17'd16873: data = 8'hf4;
      17'd16874: data = 8'h0c;
      17'd16875: data = 8'hfc;
      17'd16876: data = 8'h02;
      17'd16877: data = 8'h12;
      17'd16878: data = 8'h13;
      17'd16879: data = 8'h0c;
      17'd16880: data = 8'h0a;
      17'd16881: data = 8'h0e;
      17'd16882: data = 8'h0a;
      17'd16883: data = 8'h0a;
      17'd16884: data = 8'h06;
      17'd16885: data = 8'h12;
      17'd16886: data = 8'h12;
      17'd16887: data = 8'h12;
      17'd16888: data = 8'h1a;
      17'd16889: data = 8'h1a;
      17'd16890: data = 8'h1f;
      17'd16891: data = 8'h1b;
      17'd16892: data = 8'h1a;
      17'd16893: data = 8'h1a;
      17'd16894: data = 8'h1b;
      17'd16895: data = 8'h23;
      17'd16896: data = 8'h23;
      17'd16897: data = 8'h1f;
      17'd16898: data = 8'h1a;
      17'd16899: data = 8'h16;
      17'd16900: data = 8'h12;
      17'd16901: data = 8'h0c;
      17'd16902: data = 8'h0a;
      17'd16903: data = 8'h0a;
      17'd16904: data = 8'h0c;
      17'd16905: data = 8'h11;
      17'd16906: data = 8'h11;
      17'd16907: data = 8'h0d;
      17'd16908: data = 8'h11;
      17'd16909: data = 8'h0c;
      17'd16910: data = 8'hfd;
      17'd16911: data = 8'hf6;
      17'd16912: data = 8'hf5;
      17'd16913: data = 8'hf2;
      17'd16914: data = 8'hf2;
      17'd16915: data = 8'hef;
      17'd16916: data = 8'hec;
      17'd16917: data = 8'hef;
      17'd16918: data = 8'hec;
      17'd16919: data = 8'he4;
      17'd16920: data = 8'he4;
      17'd16921: data = 8'he7;
      17'd16922: data = 8'he7;
      17'd16923: data = 8'heb;
      17'd16924: data = 8'hef;
      17'd16925: data = 8'hec;
      17'd16926: data = 8'heb;
      17'd16927: data = 8'hef;
      17'd16928: data = 8'he5;
      17'd16929: data = 8'he5;
      17'd16930: data = 8'hef;
      17'd16931: data = 8'heb;
      17'd16932: data = 8'hef;
      17'd16933: data = 8'hf5;
      17'd16934: data = 8'hfa;
      17'd16935: data = 8'h00;
      17'd16936: data = 8'h06;
      17'd16937: data = 8'h09;
      17'd16938: data = 8'h06;
      17'd16939: data = 8'h0c;
      17'd16940: data = 8'h0e;
      17'd16941: data = 8'h0c;
      17'd16942: data = 8'h12;
      17'd16943: data = 8'h1a;
      17'd16944: data = 8'h16;
      17'd16945: data = 8'h19;
      17'd16946: data = 8'h13;
      17'd16947: data = 8'h15;
      17'd16948: data = 8'h23;
      17'd16949: data = 8'h24;
      17'd16950: data = 8'h27;
      17'd16951: data = 8'h35;
      17'd16952: data = 8'h34;
      17'd16953: data = 8'h29;
      17'd16954: data = 8'h23;
      17'd16955: data = 8'h26;
      17'd16956: data = 8'h27;
      17'd16957: data = 8'h22;
      17'd16958: data = 8'h1f;
      17'd16959: data = 8'h1b;
      17'd16960: data = 8'h1a;
      17'd16961: data = 8'h19;
      17'd16962: data = 8'h1b;
      17'd16963: data = 8'h1c;
      17'd16964: data = 8'h19;
      17'd16965: data = 8'h0d;
      17'd16966: data = 8'h13;
      17'd16967: data = 8'h0e;
      17'd16968: data = 8'hfc;
      17'd16969: data = 8'hfd;
      17'd16970: data = 8'h02;
      17'd16971: data = 8'hf2;
      17'd16972: data = 8'hed;
      17'd16973: data = 8'hfa;
      17'd16974: data = 8'hf5;
      17'd16975: data = 8'he2;
      17'd16976: data = 8'he3;
      17'd16977: data = 8'heb;
      17'd16978: data = 8'he9;
      17'd16979: data = 8'hec;
      17'd16980: data = 8'he4;
      17'd16981: data = 8'hdc;
      17'd16982: data = 8'he2;
      17'd16983: data = 8'hdc;
      17'd16984: data = 8'hd6;
      17'd16985: data = 8'hdc;
      17'd16986: data = 8'hd8;
      17'd16987: data = 8'hd3;
      17'd16988: data = 8'hdb;
      17'd16989: data = 8'hdc;
      17'd16990: data = 8'he2;
      17'd16991: data = 8'hec;
      17'd16992: data = 8'he9;
      17'd16993: data = 8'he5;
      17'd16994: data = 8'he7;
      17'd16995: data = 8'he4;
      17'd16996: data = 8'he9;
      17'd16997: data = 8'hed;
      17'd16998: data = 8'he7;
      17'd16999: data = 8'he5;
      17'd17000: data = 8'hef;
      17'd17001: data = 8'hef;
      17'd17002: data = 8'hf1;
      17'd17003: data = 8'hf9;
      17'd17004: data = 8'hf5;
      17'd17005: data = 8'hf2;
      17'd17006: data = 8'hfa;
      17'd17007: data = 8'hfa;
      17'd17008: data = 8'hfd;
      17'd17009: data = 8'h01;
      17'd17010: data = 8'hf6;
      17'd17011: data = 8'hf4;
      17'd17012: data = 8'hf6;
      17'd17013: data = 8'hf2;
      17'd17014: data = 8'hf4;
      17'd17015: data = 8'hf6;
      17'd17016: data = 8'hed;
      17'd17017: data = 8'heb;
      17'd17018: data = 8'hfa;
      17'd17019: data = 8'hfa;
      17'd17020: data = 8'hf4;
      17'd17021: data = 8'hf6;
      17'd17022: data = 8'hf4;
      17'd17023: data = 8'he9;
      17'd17024: data = 8'he9;
      17'd17025: data = 8'he9;
      17'd17026: data = 8'heb;
      17'd17027: data = 8'hec;
      17'd17028: data = 8'he5;
      17'd17029: data = 8'he3;
      17'd17030: data = 8'he7;
      17'd17031: data = 8'he9;
      17'd17032: data = 8'he4;
      17'd17033: data = 8'he7;
      17'd17034: data = 8'he9;
      17'd17035: data = 8'he7;
      17'd17036: data = 8'he9;
      17'd17037: data = 8'hed;
      17'd17038: data = 8'hed;
      17'd17039: data = 8'he9;
      17'd17040: data = 8'he9;
      17'd17041: data = 8'heb;
      17'd17042: data = 8'heb;
      17'd17043: data = 8'he7;
      17'd17044: data = 8'hec;
      17'd17045: data = 8'hf4;
      17'd17046: data = 8'hf4;
      17'd17047: data = 8'hf6;
      17'd17048: data = 8'hfe;
      17'd17049: data = 8'h04;
      17'd17050: data = 8'h00;
      17'd17051: data = 8'h01;
      17'd17052: data = 8'h06;
      17'd17053: data = 8'h00;
      17'd17054: data = 8'h00;
      17'd17055: data = 8'h09;
      17'd17056: data = 8'h0d;
      17'd17057: data = 8'h09;
      17'd17058: data = 8'h0c;
      17'd17059: data = 8'h12;
      17'd17060: data = 8'h0a;
      17'd17061: data = 8'h06;
      17'd17062: data = 8'h12;
      17'd17063: data = 8'h15;
      17'd17064: data = 8'h13;
      17'd17065: data = 8'h16;
      17'd17066: data = 8'h16;
      17'd17067: data = 8'h13;
      17'd17068: data = 8'h1f;
      17'd17069: data = 8'h1b;
      17'd17070: data = 8'h09;
      17'd17071: data = 8'h11;
      17'd17072: data = 8'h13;
      17'd17073: data = 8'h04;
      17'd17074: data = 8'h04;
      17'd17075: data = 8'h0a;
      17'd17076: data = 8'h11;
      17'd17077: data = 8'h13;
      17'd17078: data = 8'h0c;
      17'd17079: data = 8'h0a;
      17'd17080: data = 8'h0d;
      17'd17081: data = 8'h0c;
      17'd17082: data = 8'hfa;
      17'd17083: data = 8'h00;
      17'd17084: data = 8'h19;
      17'd17085: data = 8'h06;
      17'd17086: data = 8'hf5;
      17'd17087: data = 8'h0a;
      17'd17088: data = 8'h0e;
      17'd17089: data = 8'hf9;
      17'd17090: data = 8'hf5;
      17'd17091: data = 8'h02;
      17'd17092: data = 8'h05;
      17'd17093: data = 8'hf9;
      17'd17094: data = 8'hfe;
      17'd17095: data = 8'h09;
      17'd17096: data = 8'h05;
      17'd17097: data = 8'h06;
      17'd17098: data = 8'h0c;
      17'd17099: data = 8'h0a;
      17'd17100: data = 8'h05;
      17'd17101: data = 8'h06;
      17'd17102: data = 8'hfe;
      17'd17103: data = 8'hfd;
      17'd17104: data = 8'h01;
      17'd17105: data = 8'h0e;
      17'd17106: data = 8'h16;
      17'd17107: data = 8'h16;
      17'd17108: data = 8'h1e;
      17'd17109: data = 8'h26;
      17'd17110: data = 8'h1b;
      17'd17111: data = 8'h12;
      17'd17112: data = 8'h1b;
      17'd17113: data = 8'h23;
      17'd17114: data = 8'h1c;
      17'd17115: data = 8'h1a;
      17'd17116: data = 8'h24;
      17'd17117: data = 8'h29;
      17'd17118: data = 8'h1f;
      17'd17119: data = 8'h1c;
      17'd17120: data = 8'h23;
      17'd17121: data = 8'h2b;
      17'd17122: data = 8'h22;
      17'd17123: data = 8'h1e;
      17'd17124: data = 8'h2b;
      17'd17125: data = 8'h29;
      17'd17126: data = 8'h22;
      17'd17127: data = 8'h22;
      17'd17128: data = 8'h24;
      17'd17129: data = 8'h1b;
      17'd17130: data = 8'h0e;
      17'd17131: data = 8'h0a;
      17'd17132: data = 8'h0c;
      17'd17133: data = 8'h0d;
      17'd17134: data = 8'h0a;
      17'd17135: data = 8'h0c;
      17'd17136: data = 8'h0c;
      17'd17137: data = 8'h0a;
      17'd17138: data = 8'h02;
      17'd17139: data = 8'hfd;
      17'd17140: data = 8'hf9;
      17'd17141: data = 8'hf4;
      17'd17142: data = 8'hf2;
      17'd17143: data = 8'heb;
      17'd17144: data = 8'he9;
      17'd17145: data = 8'hed;
      17'd17146: data = 8'he9;
      17'd17147: data = 8'he3;
      17'd17148: data = 8'he4;
      17'd17149: data = 8'he4;
      17'd17150: data = 8'he3;
      17'd17151: data = 8'hde;
      17'd17152: data = 8'hdc;
      17'd17153: data = 8'he4;
      17'd17154: data = 8'he4;
      17'd17155: data = 8'hde;
      17'd17156: data = 8'he4;
      17'd17157: data = 8'he7;
      17'd17158: data = 8'hde;
      17'd17159: data = 8'hda;
      17'd17160: data = 8'he4;
      17'd17161: data = 8'he7;
      17'd17162: data = 8'heb;
      17'd17163: data = 8'hf2;
      17'd17164: data = 8'hf5;
      17'd17165: data = 8'hfe;
      17'd17166: data = 8'h02;
      17'd17167: data = 8'hfe;
      17'd17168: data = 8'h02;
      17'd17169: data = 8'h0a;
      17'd17170: data = 8'h01;
      17'd17171: data = 8'h02;
      17'd17172: data = 8'h0c;
      17'd17173: data = 8'h0c;
      17'd17174: data = 8'h0d;
      17'd17175: data = 8'h13;
      17'd17176: data = 8'h1a;
      17'd17177: data = 8'h1e;
      17'd17178: data = 8'h1c;
      17'd17179: data = 8'h1a;
      17'd17180: data = 8'h1f;
      17'd17181: data = 8'h1f;
      17'd17182: data = 8'h1c;
      17'd17183: data = 8'h1f;
      17'd17184: data = 8'h24;
      17'd17185: data = 8'h1c;
      17'd17186: data = 8'h1b;
      17'd17187: data = 8'h1b;
      17'd17188: data = 8'h16;
      17'd17189: data = 8'h13;
      17'd17190: data = 8'h0e;
      17'd17191: data = 8'h0d;
      17'd17192: data = 8'h16;
      17'd17193: data = 8'h11;
      17'd17194: data = 8'h0c;
      17'd17195: data = 8'h0e;
      17'd17196: data = 8'h09;
      17'd17197: data = 8'h01;
      17'd17198: data = 8'h00;
      17'd17199: data = 8'hfd;
      17'd17200: data = 8'hf6;
      17'd17201: data = 8'hf5;
      17'd17202: data = 8'hf1;
      17'd17203: data = 8'hed;
      17'd17204: data = 8'hf1;
      17'd17205: data = 8'hec;
      17'd17206: data = 8'he5;
      17'd17207: data = 8'he7;
      17'd17208: data = 8'he4;
      17'd17209: data = 8'hde;
      17'd17210: data = 8'he2;
      17'd17211: data = 8'he2;
      17'd17212: data = 8'hdc;
      17'd17213: data = 8'hde;
      17'd17214: data = 8'hde;
      17'd17215: data = 8'hde;
      17'd17216: data = 8'hdc;
      17'd17217: data = 8'hdc;
      17'd17218: data = 8'he0;
      17'd17219: data = 8'hdc;
      17'd17220: data = 8'hd8;
      17'd17221: data = 8'hde;
      17'd17222: data = 8'he4;
      17'd17223: data = 8'he4;
      17'd17224: data = 8'he4;
      17'd17225: data = 8'he4;
      17'd17226: data = 8'he4;
      17'd17227: data = 8'he4;
      17'd17228: data = 8'he5;
      17'd17229: data = 8'he7;
      17'd17230: data = 8'heb;
      17'd17231: data = 8'heb;
      17'd17232: data = 8'hef;
      17'd17233: data = 8'hed;
      17'd17234: data = 8'hf2;
      17'd17235: data = 8'hf4;
      17'd17236: data = 8'hef;
      17'd17237: data = 8'hf2;
      17'd17238: data = 8'hf4;
      17'd17239: data = 8'hf2;
      17'd17240: data = 8'hf4;
      17'd17241: data = 8'hf4;
      17'd17242: data = 8'hf5;
      17'd17243: data = 8'hf6;
      17'd17244: data = 8'hf9;
      17'd17245: data = 8'hf6;
      17'd17246: data = 8'hf5;
      17'd17247: data = 8'hfa;
      17'd17248: data = 8'hf6;
      17'd17249: data = 8'hf5;
      17'd17250: data = 8'hf9;
      17'd17251: data = 8'hfa;
      17'd17252: data = 8'hf5;
      17'd17253: data = 8'hf4;
      17'd17254: data = 8'hf9;
      17'd17255: data = 8'hf5;
      17'd17256: data = 8'hf1;
      17'd17257: data = 8'hf2;
      17'd17258: data = 8'hf4;
      17'd17259: data = 8'hf2;
      17'd17260: data = 8'hf2;
      17'd17261: data = 8'hf6;
      17'd17262: data = 8'hf5;
      17'd17263: data = 8'hf4;
      17'd17264: data = 8'hf5;
      17'd17265: data = 8'hf6;
      17'd17266: data = 8'hf5;
      17'd17267: data = 8'hf2;
      17'd17268: data = 8'hf4;
      17'd17269: data = 8'hf6;
      17'd17270: data = 8'hf4;
      17'd17271: data = 8'hef;
      17'd17272: data = 8'hf4;
      17'd17273: data = 8'hfd;
      17'd17274: data = 8'hfe;
      17'd17275: data = 8'hf9;
      17'd17276: data = 8'h01;
      17'd17277: data = 8'h00;
      17'd17278: data = 8'h00;
      17'd17279: data = 8'h00;
      17'd17280: data = 8'hfa;
      17'd17281: data = 8'h00;
      17'd17282: data = 8'h12;
      17'd17283: data = 8'h12;
      17'd17284: data = 8'h05;
      17'd17285: data = 8'h09;
      17'd17286: data = 8'h05;
      17'd17287: data = 8'h02;
      17'd17288: data = 8'h09;
      17'd17289: data = 8'h12;
      17'd17290: data = 8'h11;
      17'd17291: data = 8'h0d;
      17'd17292: data = 8'h13;
      17'd17293: data = 8'h11;
      17'd17294: data = 8'h0e;
      17'd17295: data = 8'h13;
      17'd17296: data = 8'h13;
      17'd17297: data = 8'h15;
      17'd17298: data = 8'h15;
      17'd17299: data = 8'h0e;
      17'd17300: data = 8'h0c;
      17'd17301: data = 8'h09;
      17'd17302: data = 8'h0a;
      17'd17303: data = 8'h15;
      17'd17304: data = 8'h11;
      17'd17305: data = 8'h09;
      17'd17306: data = 8'h09;
      17'd17307: data = 8'h09;
      17'd17308: data = 8'h05;
      17'd17309: data = 8'h0d;
      17'd17310: data = 8'h0e;
      17'd17311: data = 8'h0c;
      17'd17312: data = 8'h0c;
      17'd17313: data = 8'h15;
      17'd17314: data = 8'h13;
      17'd17315: data = 8'h02;
      17'd17316: data = 8'hfa;
      17'd17317: data = 8'h04;
      17'd17318: data = 8'h06;
      17'd17319: data = 8'h00;
      17'd17320: data = 8'h05;
      17'd17321: data = 8'h09;
      17'd17322: data = 8'h0a;
      17'd17323: data = 8'h0a;
      17'd17324: data = 8'h06;
      17'd17325: data = 8'h02;
      17'd17326: data = 8'h01;
      17'd17327: data = 8'h0a;
      17'd17328: data = 8'h0c;
      17'd17329: data = 8'h05;
      17'd17330: data = 8'h05;
      17'd17331: data = 8'h0a;
      17'd17332: data = 8'h09;
      17'd17333: data = 8'h04;
      17'd17334: data = 8'h0a;
      17'd17335: data = 8'h0a;
      17'd17336: data = 8'h04;
      17'd17337: data = 8'h00;
      17'd17338: data = 8'h06;
      17'd17339: data = 8'h0a;
      17'd17340: data = 8'h0a;
      17'd17341: data = 8'h0d;
      17'd17342: data = 8'h13;
      17'd17343: data = 8'h16;
      17'd17344: data = 8'h15;
      17'd17345: data = 8'h12;
      17'd17346: data = 8'h06;
      17'd17347: data = 8'h0a;
      17'd17348: data = 8'h0d;
      17'd17349: data = 8'h0e;
      17'd17350: data = 8'h12;
      17'd17351: data = 8'h11;
      17'd17352: data = 8'h13;
      17'd17353: data = 8'h15;
      17'd17354: data = 8'h0e;
      17'd17355: data = 8'h0c;
      17'd17356: data = 8'h11;
      17'd17357: data = 8'h12;
      17'd17358: data = 8'h0d;
      17'd17359: data = 8'h0e;
      17'd17360: data = 8'h13;
      17'd17361: data = 8'h15;
      17'd17362: data = 8'h0e;
      17'd17363: data = 8'h09;
      17'd17364: data = 8'h0a;
      17'd17365: data = 8'h09;
      17'd17366: data = 8'h05;
      17'd17367: data = 8'h00;
      17'd17368: data = 8'h02;
      17'd17369: data = 8'h04;
      17'd17370: data = 8'h04;
      17'd17371: data = 8'h02;
      17'd17372: data = 8'h04;
      17'd17373: data = 8'h02;
      17'd17374: data = 8'hfe;
      17'd17375: data = 8'hfd;
      17'd17376: data = 8'hf6;
      17'd17377: data = 8'hf6;
      17'd17378: data = 8'hf6;
      17'd17379: data = 8'hf5;
      17'd17380: data = 8'hf6;
      17'd17381: data = 8'hf5;
      17'd17382: data = 8'hf5;
      17'd17383: data = 8'hf4;
      17'd17384: data = 8'hf1;
      17'd17385: data = 8'hef;
      17'd17386: data = 8'hef;
      17'd17387: data = 8'hed;
      17'd17388: data = 8'hf1;
      17'd17389: data = 8'hf2;
      17'd17390: data = 8'hf2;
      17'd17391: data = 8'hf1;
      17'd17392: data = 8'hef;
      17'd17393: data = 8'hed;
      17'd17394: data = 8'hec;
      17'd17395: data = 8'heb;
      17'd17396: data = 8'hec;
      17'd17397: data = 8'hf2;
      17'd17398: data = 8'hf2;
      17'd17399: data = 8'hef;
      17'd17400: data = 8'hf4;
      17'd17401: data = 8'hf9;
      17'd17402: data = 8'hf6;
      17'd17403: data = 8'hf4;
      17'd17404: data = 8'hfa;
      17'd17405: data = 8'hf9;
      17'd17406: data = 8'hf9;
      17'd17407: data = 8'hfc;
      17'd17408: data = 8'hfc;
      17'd17409: data = 8'hfe;
      17'd17410: data = 8'hfe;
      17'd17411: data = 8'h00;
      17'd17412: data = 8'hfe;
      17'd17413: data = 8'hfe;
      17'd17414: data = 8'h02;
      17'd17415: data = 8'h05;
      17'd17416: data = 8'h05;
      17'd17417: data = 8'h09;
      17'd17418: data = 8'h06;
      17'd17419: data = 8'h06;
      17'd17420: data = 8'h09;
      17'd17421: data = 8'h09;
      17'd17422: data = 8'h09;
      17'd17423: data = 8'h06;
      17'd17424: data = 8'h05;
      17'd17425: data = 8'h06;
      17'd17426: data = 8'h06;
      17'd17427: data = 8'h09;
      17'd17428: data = 8'h09;
      17'd17429: data = 8'h05;
      17'd17430: data = 8'h05;
      17'd17431: data = 8'h04;
      17'd17432: data = 8'h02;
      17'd17433: data = 8'h02;
      17'd17434: data = 8'h02;
      17'd17435: data = 8'hfe;
      17'd17436: data = 8'hfd;
      17'd17437: data = 8'h00;
      17'd17438: data = 8'hfd;
      17'd17439: data = 8'hfd;
      17'd17440: data = 8'hfd;
      17'd17441: data = 8'hfa;
      17'd17442: data = 8'hf5;
      17'd17443: data = 8'hf4;
      17'd17444: data = 8'hf4;
      17'd17445: data = 8'hf2;
      17'd17446: data = 8'hf2;
      17'd17447: data = 8'hf2;
      17'd17448: data = 8'hf2;
      17'd17449: data = 8'hf2;
      17'd17450: data = 8'hf1;
      17'd17451: data = 8'hed;
      17'd17452: data = 8'hec;
      17'd17453: data = 8'hec;
      17'd17454: data = 8'hed;
      17'd17455: data = 8'hec;
      17'd17456: data = 8'hed;
      17'd17457: data = 8'heb;
      17'd17458: data = 8'hec;
      17'd17459: data = 8'hef;
      17'd17460: data = 8'heb;
      17'd17461: data = 8'he7;
      17'd17462: data = 8'heb;
      17'd17463: data = 8'heb;
      17'd17464: data = 8'heb;
      17'd17465: data = 8'hec;
      17'd17466: data = 8'hef;
      17'd17467: data = 8'hed;
      17'd17468: data = 8'hec;
      17'd17469: data = 8'hef;
      17'd17470: data = 8'hf1;
      17'd17471: data = 8'hed;
      17'd17472: data = 8'hef;
      17'd17473: data = 8'hef;
      17'd17474: data = 8'hed;
      17'd17475: data = 8'hf2;
      17'd17476: data = 8'hf4;
      17'd17477: data = 8'hf2;
      17'd17478: data = 8'hf4;
      17'd17479: data = 8'hf4;
      17'd17480: data = 8'hf4;
      17'd17481: data = 8'hf4;
      17'd17482: data = 8'hf4;
      17'd17483: data = 8'hf4;
      17'd17484: data = 8'hf5;
      17'd17485: data = 8'hf4;
      17'd17486: data = 8'hf5;
      17'd17487: data = 8'hfa;
      17'd17488: data = 8'hfa;
      17'd17489: data = 8'hf5;
      17'd17490: data = 8'hf6;
      17'd17491: data = 8'hf9;
      17'd17492: data = 8'hfc;
      17'd17493: data = 8'hfa;
      17'd17494: data = 8'hf5;
      17'd17495: data = 8'hf9;
      17'd17496: data = 8'hfa;
      17'd17497: data = 8'hf9;
      17'd17498: data = 8'hf6;
      17'd17499: data = 8'hfa;
      17'd17500: data = 8'hfa;
      17'd17501: data = 8'hf9;
      17'd17502: data = 8'hfa;
      17'd17503: data = 8'hfc;
      17'd17504: data = 8'hfc;
      17'd17505: data = 8'hfc;
      17'd17506: data = 8'hfe;
      17'd17507: data = 8'hfd;
      17'd17508: data = 8'hfd;
      17'd17509: data = 8'h00;
      17'd17510: data = 8'h00;
      17'd17511: data = 8'hfe;
      17'd17512: data = 8'h02;
      17'd17513: data = 8'h04;
      17'd17514: data = 8'h01;
      17'd17515: data = 8'h04;
      17'd17516: data = 8'h05;
      17'd17517: data = 8'h02;
      17'd17518: data = 8'h06;
      17'd17519: data = 8'h09;
      17'd17520: data = 8'h04;
      17'd17521: data = 8'h06;
      17'd17522: data = 8'h0d;
      17'd17523: data = 8'h0c;
      17'd17524: data = 8'h05;
      17'd17525: data = 8'h09;
      17'd17526: data = 8'h0c;
      17'd17527: data = 8'h0d;
      17'd17528: data = 8'h0d;
      17'd17529: data = 8'h0c;
      17'd17530: data = 8'h0d;
      17'd17531: data = 8'h0e;
      17'd17532: data = 8'h0d;
      17'd17533: data = 8'h11;
      17'd17534: data = 8'h0e;
      17'd17535: data = 8'h0c;
      17'd17536: data = 8'h0a;
      17'd17537: data = 8'h0e;
      17'd17538: data = 8'h0d;
      17'd17539: data = 8'h0d;
      17'd17540: data = 8'h0e;
      17'd17541: data = 8'h0c;
      17'd17542: data = 8'h0d;
      17'd17543: data = 8'h11;
      17'd17544: data = 8'h0e;
      17'd17545: data = 8'h0a;
      17'd17546: data = 8'h0c;
      17'd17547: data = 8'h0e;
      17'd17548: data = 8'h11;
      17'd17549: data = 8'h0d;
      17'd17550: data = 8'h0c;
      17'd17551: data = 8'h0d;
      17'd17552: data = 8'h0c;
      17'd17553: data = 8'h0d;
      17'd17554: data = 8'h0e;
      17'd17555: data = 8'h0a;
      17'd17556: data = 8'h0a;
      17'd17557: data = 8'h0c;
      17'd17558: data = 8'h0e;
      17'd17559: data = 8'h0a;
      17'd17560: data = 8'h05;
      17'd17561: data = 8'h05;
      17'd17562: data = 8'h09;
      17'd17563: data = 8'h06;
      17'd17564: data = 8'h04;
      17'd17565: data = 8'h06;
      17'd17566: data = 8'h09;
      17'd17567: data = 8'h09;
      17'd17568: data = 8'h05;
      17'd17569: data = 8'h02;
      17'd17570: data = 8'h05;
      17'd17571: data = 8'h06;
      17'd17572: data = 8'h04;
      17'd17573: data = 8'h00;
      17'd17574: data = 8'h04;
      17'd17575: data = 8'h05;
      17'd17576: data = 8'h02;
      17'd17577: data = 8'h02;
      17'd17578: data = 8'h00;
      17'd17579: data = 8'h00;
      17'd17580: data = 8'h01;
      17'd17581: data = 8'h00;
      17'd17582: data = 8'hfd;
      17'd17583: data = 8'hfe;
      17'd17584: data = 8'h01;
      17'd17585: data = 8'hfe;
      17'd17586: data = 8'hfd;
      17'd17587: data = 8'hfe;
      17'd17588: data = 8'h02;
      17'd17589: data = 8'h02;
      17'd17590: data = 8'hfd;
      17'd17591: data = 8'hfc;
      17'd17592: data = 8'h01;
      17'd17593: data = 8'h01;
      17'd17594: data = 8'h00;
      17'd17595: data = 8'h00;
      17'd17596: data = 8'h00;
      17'd17597: data = 8'h02;
      17'd17598: data = 8'h04;
      17'd17599: data = 8'h02;
      17'd17600: data = 8'h01;
      17'd17601: data = 8'hfe;
      17'd17602: data = 8'h00;
      17'd17603: data = 8'h05;
      17'd17604: data = 8'h01;
      17'd17605: data = 8'hfe;
      17'd17606: data = 8'h04;
      17'd17607: data = 8'h04;
      17'd17608: data = 8'hfe;
      17'd17609: data = 8'h01;
      17'd17610: data = 8'h02;
      17'd17611: data = 8'h00;
      17'd17612: data = 8'h01;
      17'd17613: data = 8'h02;
      17'd17614: data = 8'h02;
      17'd17615: data = 8'h02;
      17'd17616: data = 8'h04;
      17'd17617: data = 8'h01;
      17'd17618: data = 8'hfe;
      17'd17619: data = 8'h02;
      17'd17620: data = 8'h01;
      17'd17621: data = 8'h00;
      17'd17622: data = 8'hfe;
      17'd17623: data = 8'hfd;
      17'd17624: data = 8'hfd;
      17'd17625: data = 8'h00;
      17'd17626: data = 8'hfe;
      17'd17627: data = 8'hfc;
      17'd17628: data = 8'hfa;
      17'd17629: data = 8'hf5;
      17'd17630: data = 8'hf6;
      17'd17631: data = 8'hf6;
      17'd17632: data = 8'hf5;
      17'd17633: data = 8'hf6;
      17'd17634: data = 8'hf6;
      17'd17635: data = 8'hf4;
      17'd17636: data = 8'hf2;
      17'd17637: data = 8'hf4;
      17'd17638: data = 8'hf6;
      17'd17639: data = 8'hf2;
      17'd17640: data = 8'hef;
      17'd17641: data = 8'hf5;
      17'd17642: data = 8'hf5;
      17'd17643: data = 8'hf1;
      17'd17644: data = 8'hf2;
      17'd17645: data = 8'hf4;
      17'd17646: data = 8'hf4;
      17'd17647: data = 8'hf2;
      17'd17648: data = 8'hf2;
      17'd17649: data = 8'hf2;
      17'd17650: data = 8'hf4;
      17'd17651: data = 8'hf4;
      17'd17652: data = 8'hf4;
      17'd17653: data = 8'hf5;
      17'd17654: data = 8'hf4;
      17'd17655: data = 8'hf5;
      17'd17656: data = 8'hf9;
      17'd17657: data = 8'hf6;
      17'd17658: data = 8'hf5;
      17'd17659: data = 8'hf9;
      17'd17660: data = 8'hfc;
      17'd17661: data = 8'hfc;
      17'd17662: data = 8'hfc;
      17'd17663: data = 8'hfd;
      17'd17664: data = 8'hfe;
      17'd17665: data = 8'h00;
      17'd17666: data = 8'h01;
      17'd17667: data = 8'hfe;
      17'd17668: data = 8'h01;
      17'd17669: data = 8'h01;
      17'd17670: data = 8'h01;
      17'd17671: data = 8'h02;
      17'd17672: data = 8'h04;
      17'd17673: data = 8'h04;
      17'd17674: data = 8'h04;
      17'd17675: data = 8'h02;
      17'd17676: data = 8'h04;
      17'd17677: data = 8'h05;
      17'd17678: data = 8'h06;
      17'd17679: data = 8'h06;
      17'd17680: data = 8'h04;
      17'd17681: data = 8'h05;
      17'd17682: data = 8'h06;
      17'd17683: data = 8'h09;
      17'd17684: data = 8'h06;
      17'd17685: data = 8'h05;
      17'd17686: data = 8'h05;
      17'd17687: data = 8'h05;
      17'd17688: data = 8'h04;
      17'd17689: data = 8'h05;
      17'd17690: data = 8'h09;
      17'd17691: data = 8'h05;
      17'd17692: data = 8'h02;
      17'd17693: data = 8'h05;
      17'd17694: data = 8'h06;
      17'd17695: data = 8'h04;
      17'd17696: data = 8'h01;
      17'd17697: data = 8'h01;
      17'd17698: data = 8'h01;
      17'd17699: data = 8'h01;
      17'd17700: data = 8'h01;
      17'd17701: data = 8'h02;
      17'd17702: data = 8'h01;
      17'd17703: data = 8'h00;
      17'd17704: data = 8'hfd;
      17'd17705: data = 8'hfd;
      17'd17706: data = 8'h00;
      17'd17707: data = 8'h00;
      17'd17708: data = 8'hfd;
      17'd17709: data = 8'hfd;
      17'd17710: data = 8'hfd;
      17'd17711: data = 8'hfd;
      17'd17712: data = 8'h00;
      17'd17713: data = 8'hfa;
      17'd17714: data = 8'hf6;
      17'd17715: data = 8'hfa;
      17'd17716: data = 8'hf9;
      17'd17717: data = 8'hf5;
      17'd17718: data = 8'hfa;
      17'd17719: data = 8'hf9;
      17'd17720: data = 8'hf5;
      17'd17721: data = 8'hf9;
      17'd17722: data = 8'hfc;
      17'd17723: data = 8'hf5;
      17'd17724: data = 8'hf4;
      17'd17725: data = 8'hfa;
      17'd17726: data = 8'hf6;
      17'd17727: data = 8'hf5;
      17'd17728: data = 8'hf5;
      17'd17729: data = 8'hf6;
      17'd17730: data = 8'hf5;
      17'd17731: data = 8'hf6;
      17'd17732: data = 8'hf6;
      17'd17733: data = 8'hf2;
      17'd17734: data = 8'hf2;
      17'd17735: data = 8'hf6;
      17'd17736: data = 8'hf6;
      17'd17737: data = 8'hf5;
      17'd17738: data = 8'hf6;
      17'd17739: data = 8'hf5;
      17'd17740: data = 8'hf6;
      17'd17741: data = 8'hf6;
      17'd17742: data = 8'hf6;
      17'd17743: data = 8'hf5;
      17'd17744: data = 8'hef;
      17'd17745: data = 8'hf2;
      17'd17746: data = 8'hf5;
      17'd17747: data = 8'hf6;
      17'd17748: data = 8'hf5;
      17'd17749: data = 8'hf5;
      17'd17750: data = 8'hf6;
      17'd17751: data = 8'hf5;
      17'd17752: data = 8'hf5;
      17'd17753: data = 8'hf6;
      17'd17754: data = 8'hf4;
      17'd17755: data = 8'hf5;
      17'd17756: data = 8'hf6;
      17'd17757: data = 8'hf5;
      17'd17758: data = 8'hf6;
      17'd17759: data = 8'hf5;
      17'd17760: data = 8'hf5;
      17'd17761: data = 8'hfa;
      17'd17762: data = 8'hfc;
      17'd17763: data = 8'hfa;
      17'd17764: data = 8'hfa;
      17'd17765: data = 8'hfc;
      17'd17766: data = 8'hfc;
      17'd17767: data = 8'hfe;
      17'd17768: data = 8'hfe;
      17'd17769: data = 8'hfe;
      17'd17770: data = 8'h00;
      17'd17771: data = 8'h02;
      17'd17772: data = 8'h01;
      17'd17773: data = 8'hfc;
      17'd17774: data = 8'h00;
      17'd17775: data = 8'h04;
      17'd17776: data = 8'h02;
      17'd17777: data = 8'h02;
      17'd17778: data = 8'h04;
      17'd17779: data = 8'h09;
      17'd17780: data = 8'h0a;
      17'd17781: data = 8'h05;
      17'd17782: data = 8'h05;
      17'd17783: data = 8'h0d;
      17'd17784: data = 8'h11;
      17'd17785: data = 8'h0a;
      17'd17786: data = 8'h0a;
      17'd17787: data = 8'h0d;
      17'd17788: data = 8'h0c;
      17'd17789: data = 8'h0c;
      17'd17790: data = 8'h0d;
      17'd17791: data = 8'h0d;
      17'd17792: data = 8'h0e;
      17'd17793: data = 8'h0e;
      17'd17794: data = 8'h0e;
      17'd17795: data = 8'h11;
      17'd17796: data = 8'h12;
      17'd17797: data = 8'h11;
      17'd17798: data = 8'h0e;
      17'd17799: data = 8'h12;
      17'd17800: data = 8'h12;
      17'd17801: data = 8'h0d;
      17'd17802: data = 8'h0d;
      17'd17803: data = 8'h0e;
      17'd17804: data = 8'h0e;
      17'd17805: data = 8'h0d;
      17'd17806: data = 8'h0c;
      17'd17807: data = 8'h0a;
      17'd17808: data = 8'h0c;
      17'd17809: data = 8'h0d;
      17'd17810: data = 8'h0c;
      17'd17811: data = 8'h0a;
      17'd17812: data = 8'h09;
      17'd17813: data = 8'h09;
      17'd17814: data = 8'h09;
      17'd17815: data = 8'h05;
      17'd17816: data = 8'h04;
      17'd17817: data = 8'h04;
      17'd17818: data = 8'h05;
      17'd17819: data = 8'h02;
      17'd17820: data = 8'h00;
      17'd17821: data = 8'h00;
      17'd17822: data = 8'h00;
      17'd17823: data = 8'h00;
      17'd17824: data = 8'h05;
      17'd17825: data = 8'h01;
      17'd17826: data = 8'hfd;
      17'd17827: data = 8'h00;
      17'd17828: data = 8'h01;
      17'd17829: data = 8'hfa;
      17'd17830: data = 8'hf9;
      17'd17831: data = 8'hfd;
      17'd17832: data = 8'hfd;
      17'd17833: data = 8'h01;
      17'd17834: data = 8'h00;
      17'd17835: data = 8'hfa;
      17'd17836: data = 8'hfd;
      17'd17837: data = 8'h01;
      17'd17838: data = 8'h04;
      17'd17839: data = 8'hfe;
      17'd17840: data = 8'h00;
      17'd17841: data = 8'h04;
      17'd17842: data = 8'h02;
      17'd17843: data = 8'h04;
      17'd17844: data = 8'h04;
      17'd17845: data = 8'h04;
      17'd17846: data = 8'h05;
      17'd17847: data = 8'h09;
      17'd17848: data = 8'h02;
      17'd17849: data = 8'h05;
      17'd17850: data = 8'h0c;
      17'd17851: data = 8'h09;
      17'd17852: data = 8'h0c;
      17'd17853: data = 8'h0d;
      17'd17854: data = 8'h0c;
      17'd17855: data = 8'h0d;
      17'd17856: data = 8'h12;
      17'd17857: data = 8'h0e;
      17'd17858: data = 8'h0a;
      17'd17859: data = 8'h0c;
      17'd17860: data = 8'h0e;
      17'd17861: data = 8'h0c;
      17'd17862: data = 8'h0a;
      17'd17863: data = 8'h0c;
      17'd17864: data = 8'h09;
      17'd17865: data = 8'h09;
      17'd17866: data = 8'h0c;
      17'd17867: data = 8'h09;
      17'd17868: data = 8'h06;
      17'd17869: data = 8'h0a;
      17'd17870: data = 8'h05;
      17'd17871: data = 8'h04;
      17'd17872: data = 8'h05;
      17'd17873: data = 8'h02;
      17'd17874: data = 8'h00;
      17'd17875: data = 8'h00;
      17'd17876: data = 8'hfe;
      17'd17877: data = 8'hfc;
      17'd17878: data = 8'hfc;
      17'd17879: data = 8'hfc;
      17'd17880: data = 8'hf9;
      17'd17881: data = 8'hf6;
      17'd17882: data = 8'hfa;
      17'd17883: data = 8'hf9;
      17'd17884: data = 8'hf6;
      17'd17885: data = 8'hf6;
      17'd17886: data = 8'hf5;
      17'd17887: data = 8'hf4;
      17'd17888: data = 8'hf6;
      17'd17889: data = 8'hf4;
      17'd17890: data = 8'hef;
      17'd17891: data = 8'hf4;
      17'd17892: data = 8'hf4;
      17'd17893: data = 8'hf4;
      17'd17894: data = 8'hf2;
      17'd17895: data = 8'hf4;
      17'd17896: data = 8'hf6;
      17'd17897: data = 8'hf9;
      17'd17898: data = 8'hfa;
      17'd17899: data = 8'hf6;
      17'd17900: data = 8'hf6;
      17'd17901: data = 8'hf9;
      17'd17902: data = 8'hfc;
      17'd17903: data = 8'hfa;
      17'd17904: data = 8'hf9;
      17'd17905: data = 8'hf9;
      17'd17906: data = 8'hfc;
      17'd17907: data = 8'hfc;
      17'd17908: data = 8'hfc;
      17'd17909: data = 8'hfe;
      17'd17910: data = 8'hfe;
      17'd17911: data = 8'h00;
      17'd17912: data = 8'h02;
      17'd17913: data = 8'h02;
      17'd17914: data = 8'h00;
      17'd17915: data = 8'h01;
      17'd17916: data = 8'h04;
      17'd17917: data = 8'h02;
      17'd17918: data = 8'h00;
      17'd17919: data = 8'h01;
      17'd17920: data = 8'h04;
      17'd17921: data = 8'h02;
      17'd17922: data = 8'h01;
      17'd17923: data = 8'h01;
      17'd17924: data = 8'h01;
      17'd17925: data = 8'h01;
      17'd17926: data = 8'h01;
      17'd17927: data = 8'h00;
      17'd17928: data = 8'h01;
      17'd17929: data = 8'h02;
      17'd17930: data = 8'h02;
      17'd17931: data = 8'h01;
      17'd17932: data = 8'hfe;
      17'd17933: data = 8'hfd;
      17'd17934: data = 8'h00;
      17'd17935: data = 8'h00;
      17'd17936: data = 8'hfe;
      17'd17937: data = 8'h00;
      17'd17938: data = 8'hfe;
      17'd17939: data = 8'hfc;
      17'd17940: data = 8'hfd;
      17'd17941: data = 8'hfc;
      17'd17942: data = 8'hf9;
      17'd17943: data = 8'hf6;
      17'd17944: data = 8'hfa;
      17'd17945: data = 8'hfc;
      17'd17946: data = 8'hfc;
      17'd17947: data = 8'hfa;
      17'd17948: data = 8'hfa;
      17'd17949: data = 8'hfa;
      17'd17950: data = 8'hfa;
      17'd17951: data = 8'hfa;
      17'd17952: data = 8'hfa;
      17'd17953: data = 8'hf9;
      17'd17954: data = 8'hf5;
      17'd17955: data = 8'hf9;
      17'd17956: data = 8'hf9;
      17'd17957: data = 8'hfa;
      17'd17958: data = 8'hfa;
      17'd17959: data = 8'hf5;
      17'd17960: data = 8'hf6;
      17'd17961: data = 8'hf9;
      17'd17962: data = 8'hf9;
      17'd17963: data = 8'hf9;
      17'd17964: data = 8'hf5;
      17'd17965: data = 8'hf6;
      17'd17966: data = 8'hf9;
      17'd17967: data = 8'hf4;
      17'd17968: data = 8'hf5;
      17'd17969: data = 8'hf5;
      17'd17970: data = 8'hf1;
      17'd17971: data = 8'hf1;
      17'd17972: data = 8'hf4;
      17'd17973: data = 8'hf2;
      17'd17974: data = 8'hef;
      17'd17975: data = 8'hf2;
      17'd17976: data = 8'hf2;
      17'd17977: data = 8'hf2;
      17'd17978: data = 8'hf4;
      17'd17979: data = 8'hf4;
      17'd17980: data = 8'hf4;
      17'd17981: data = 8'hf2;
      17'd17982: data = 8'hf1;
      17'd17983: data = 8'hf1;
      17'd17984: data = 8'hef;
      17'd17985: data = 8'hef;
      17'd17986: data = 8'hef;
      17'd17987: data = 8'hed;
      17'd17988: data = 8'hec;
      17'd17989: data = 8'hed;
      17'd17990: data = 8'hef;
      17'd17991: data = 8'hec;
      17'd17992: data = 8'hed;
      17'd17993: data = 8'hf1;
      17'd17994: data = 8'hf1;
      17'd17995: data = 8'hef;
      17'd17996: data = 8'hf2;
      17'd17997: data = 8'hf1;
      17'd17998: data = 8'hed;
      17'd17999: data = 8'hf1;
      17'd18000: data = 8'hf4;
      17'd18001: data = 8'hf4;
      17'd18002: data = 8'hf2;
      17'd18003: data = 8'hf2;
      17'd18004: data = 8'hf5;
      17'd18005: data = 8'hf5;
      17'd18006: data = 8'hf6;
      17'd18007: data = 8'hfc;
      17'd18008: data = 8'hfa;
      17'd18009: data = 8'hf9;
      17'd18010: data = 8'hfa;
      17'd18011: data = 8'h00;
      17'd18012: data = 8'h02;
      17'd18013: data = 8'h00;
      17'd18014: data = 8'h00;
      17'd18015: data = 8'h04;
      17'd18016: data = 8'h04;
      17'd18017: data = 8'h01;
      17'd18018: data = 8'h05;
      17'd18019: data = 8'h06;
      17'd18020: data = 8'h06;
      17'd18021: data = 8'h0c;
      17'd18022: data = 8'h0a;
      17'd18023: data = 8'h0d;
      17'd18024: data = 8'h0a;
      17'd18025: data = 8'h0c;
      17'd18026: data = 8'h0e;
      17'd18027: data = 8'h11;
      17'd18028: data = 8'h11;
      17'd18029: data = 8'h11;
      17'd18030: data = 8'h0e;
      17'd18031: data = 8'h11;
      17'd18032: data = 8'h15;
      17'd18033: data = 8'h15;
      17'd18034: data = 8'h11;
      17'd18035: data = 8'h0e;
      17'd18036: data = 8'h12;
      17'd18037: data = 8'h12;
      17'd18038: data = 8'h0e;
      17'd18039: data = 8'h0d;
      17'd18040: data = 8'h11;
      17'd18041: data = 8'h11;
      17'd18042: data = 8'h12;
      17'd18043: data = 8'h0e;
      17'd18044: data = 8'h0e;
      17'd18045: data = 8'h0e;
      17'd18046: data = 8'h0d;
      17'd18047: data = 8'h0e;
      17'd18048: data = 8'h0c;
      17'd18049: data = 8'h09;
      17'd18050: data = 8'h0a;
      17'd18051: data = 8'h0d;
      17'd18052: data = 8'h09;
      17'd18053: data = 8'h09;
      17'd18054: data = 8'h0c;
      17'd18055: data = 8'h05;
      17'd18056: data = 8'h04;
      17'd18057: data = 8'h09;
      17'd18058: data = 8'h06;
      17'd18059: data = 8'h06;
      17'd18060: data = 8'h05;
      17'd18061: data = 8'h05;
      17'd18062: data = 8'h04;
      17'd18063: data = 8'h04;
      17'd18064: data = 8'h04;
      17'd18065: data = 8'h02;
      17'd18066: data = 8'h04;
      17'd18067: data = 8'h01;
      17'd18068: data = 8'h01;
      17'd18069: data = 8'h02;
      17'd18070: data = 8'h00;
      17'd18071: data = 8'h00;
      17'd18072: data = 8'h02;
      17'd18073: data = 8'h00;
      17'd18074: data = 8'h05;
      17'd18075: data = 8'h09;
      17'd18076: data = 8'h09;
      17'd18077: data = 8'h09;
      17'd18078: data = 8'h05;
      17'd18079: data = 8'h04;
      17'd18080: data = 8'h04;
      17'd18081: data = 8'h05;
      17'd18082: data = 8'h05;
      17'd18083: data = 8'h05;
      17'd18084: data = 8'h06;
      17'd18085: data = 8'h0a;
      17'd18086: data = 8'h0d;
      17'd18087: data = 8'h0d;
      17'd18088: data = 8'h0c;
      17'd18089: data = 8'h0a;
      17'd18090: data = 8'h0d;
      17'd18091: data = 8'h11;
      17'd18092: data = 8'h0d;
      17'd18093: data = 8'h0a;
      17'd18094: data = 8'h0e;
      17'd18095: data = 8'h11;
      17'd18096: data = 8'h0d;
      17'd18097: data = 8'h0d;
      17'd18098: data = 8'h0d;
      17'd18099: data = 8'h09;
      17'd18100: data = 8'h0c;
      17'd18101: data = 8'h0e;
      17'd18102: data = 8'h0a;
      17'd18103: data = 8'h0c;
      17'd18104: data = 8'h0e;
      17'd18105: data = 8'h11;
      17'd18106: data = 8'h0a;
      17'd18107: data = 8'h05;
      17'd18108: data = 8'h06;
      17'd18109: data = 8'h0a;
      17'd18110: data = 8'h05;
      17'd18111: data = 8'h01;
      17'd18112: data = 8'h02;
      17'd18113: data = 8'hfe;
      17'd18114: data = 8'hfe;
      17'd18115: data = 8'hfe;
      17'd18116: data = 8'hfc;
      17'd18117: data = 8'hfa;
      17'd18118: data = 8'hfa;
      17'd18119: data = 8'hfa;
      17'd18120: data = 8'hf6;
      17'd18121: data = 8'hf6;
      17'd18122: data = 8'hf4;
      17'd18123: data = 8'hf5;
      17'd18124: data = 8'hf9;
      17'd18125: data = 8'hf4;
      17'd18126: data = 8'hf4;
      17'd18127: data = 8'hf4;
      17'd18128: data = 8'hf1;
      17'd18129: data = 8'hef;
      17'd18130: data = 8'hf1;
      17'd18131: data = 8'hf1;
      17'd18132: data = 8'hf1;
      17'd18133: data = 8'hef;
      17'd18134: data = 8'hef;
      17'd18135: data = 8'hef;
      17'd18136: data = 8'hf1;
      17'd18137: data = 8'hf2;
      17'd18138: data = 8'hf2;
      17'd18139: data = 8'hf4;
      17'd18140: data = 8'hf4;
      17'd18141: data = 8'hf2;
      17'd18142: data = 8'hf2;
      17'd18143: data = 8'hf2;
      17'd18144: data = 8'hf4;
      17'd18145: data = 8'hf6;
      17'd18146: data = 8'hf6;
      17'd18147: data = 8'hf6;
      17'd18148: data = 8'hf5;
      17'd18149: data = 8'hf6;
      17'd18150: data = 8'hfa;
      17'd18151: data = 8'hf9;
      17'd18152: data = 8'hf9;
      17'd18153: data = 8'hfa;
      17'd18154: data = 8'hfa;
      17'd18155: data = 8'hfa;
      17'd18156: data = 8'h01;
      17'd18157: data = 8'h00;
      17'd18158: data = 8'hfa;
      17'd18159: data = 8'hfd;
      17'd18160: data = 8'hfd;
      17'd18161: data = 8'hfd;
      17'd18162: data = 8'hfe;
      17'd18163: data = 8'hf9;
      17'd18164: data = 8'hfa;
      17'd18165: data = 8'hfd;
      17'd18166: data = 8'hfc;
      17'd18167: data = 8'hfa;
      17'd18168: data = 8'hfc;
      17'd18169: data = 8'h00;
      17'd18170: data = 8'h02;
      17'd18171: data = 8'hfe;
      17'd18172: data = 8'hfa;
      17'd18173: data = 8'hfc;
      17'd18174: data = 8'hfe;
      17'd18175: data = 8'h00;
      17'd18176: data = 8'hfc;
      17'd18177: data = 8'hf6;
      17'd18178: data = 8'hf9;
      17'd18179: data = 8'hfa;
      17'd18180: data = 8'hfc;
      17'd18181: data = 8'hf6;
      17'd18182: data = 8'hf5;
      17'd18183: data = 8'hf5;
      17'd18184: data = 8'hf9;
      17'd18185: data = 8'hfa;
      17'd18186: data = 8'hf6;
      17'd18187: data = 8'hfa;
      17'd18188: data = 8'hfc;
      17'd18189: data = 8'hfa;
      17'd18190: data = 8'hf6;
      17'd18191: data = 8'hf9;
      17'd18192: data = 8'hfa;
      17'd18193: data = 8'hf6;
      17'd18194: data = 8'hf5;
      17'd18195: data = 8'hf5;
      17'd18196: data = 8'hf5;
      17'd18197: data = 8'hf2;
      17'd18198: data = 8'hf6;
      17'd18199: data = 8'hf9;
      17'd18200: data = 8'hf4;
      17'd18201: data = 8'hf5;
      17'd18202: data = 8'hf9;
      17'd18203: data = 8'hf6;
      17'd18204: data = 8'hf5;
      17'd18205: data = 8'hf5;
      17'd18206: data = 8'hf4;
      17'd18207: data = 8'hf4;
      17'd18208: data = 8'hf4;
      17'd18209: data = 8'hf2;
      17'd18210: data = 8'hf1;
      17'd18211: data = 8'hef;
      17'd18212: data = 8'hed;
      17'd18213: data = 8'hf2;
      17'd18214: data = 8'hf2;
      17'd18215: data = 8'hec;
      17'd18216: data = 8'hef;
      17'd18217: data = 8'hf1;
      17'd18218: data = 8'hed;
      17'd18219: data = 8'hef;
      17'd18220: data = 8'hed;
      17'd18221: data = 8'hef;
      17'd18222: data = 8'hef;
      17'd18223: data = 8'hef;
      17'd18224: data = 8'hed;
      17'd18225: data = 8'hec;
      17'd18226: data = 8'hef;
      17'd18227: data = 8'hef;
      17'd18228: data = 8'hf1;
      17'd18229: data = 8'hf4;
      17'd18230: data = 8'hf4;
      17'd18231: data = 8'hf1;
      17'd18232: data = 8'hf1;
      17'd18233: data = 8'hf1;
      17'd18234: data = 8'hf5;
      17'd18235: data = 8'hf4;
      17'd18236: data = 8'hf2;
      17'd18237: data = 8'hf4;
      17'd18238: data = 8'hf2;
      17'd18239: data = 8'hf4;
      17'd18240: data = 8'hf5;
      17'd18241: data = 8'hfc;
      17'd18242: data = 8'hfd;
      17'd18243: data = 8'hfc;
      17'd18244: data = 8'hfd;
      17'd18245: data = 8'h00;
      17'd18246: data = 8'hfe;
      17'd18247: data = 8'h00;
      17'd18248: data = 8'h01;
      17'd18249: data = 8'h01;
      17'd18250: data = 8'h02;
      17'd18251: data = 8'h06;
      17'd18252: data = 8'h01;
      17'd18253: data = 8'h01;
      17'd18254: data = 8'h0a;
      17'd18255: data = 8'h0c;
      17'd18256: data = 8'h0a;
      17'd18257: data = 8'h0c;
      17'd18258: data = 8'h0d;
      17'd18259: data = 8'h0c;
      17'd18260: data = 8'h0d;
      17'd18261: data = 8'h15;
      17'd18262: data = 8'h12;
      17'd18263: data = 8'h0e;
      17'd18264: data = 8'h11;
      17'd18265: data = 8'h12;
      17'd18266: data = 8'h12;
      17'd18267: data = 8'h11;
      17'd18268: data = 8'h0e;
      17'd18269: data = 8'h13;
      17'd18270: data = 8'h12;
      17'd18271: data = 8'h13;
      17'd18272: data = 8'h16;
      17'd18273: data = 8'h16;
      17'd18274: data = 8'h13;
      17'd18275: data = 8'h13;
      17'd18276: data = 8'h13;
      17'd18277: data = 8'h13;
      17'd18278: data = 8'h13;
      17'd18279: data = 8'h12;
      17'd18280: data = 8'h12;
      17'd18281: data = 8'h0e;
      17'd18282: data = 8'h0e;
      17'd18283: data = 8'h0e;
      17'd18284: data = 8'h09;
      17'd18285: data = 8'h0e;
      17'd18286: data = 8'h12;
      17'd18287: data = 8'h11;
      17'd18288: data = 8'h11;
      17'd18289: data = 8'h0d;
      17'd18290: data = 8'h0d;
      17'd18291: data = 8'h11;
      17'd18292: data = 8'h0c;
      17'd18293: data = 8'h0a;
      17'd18294: data = 8'h0d;
      17'd18295: data = 8'h09;
      17'd18296: data = 8'h0a;
      17'd18297: data = 8'h0c;
      17'd18298: data = 8'h09;
      17'd18299: data = 8'h06;
      17'd18300: data = 8'h0a;
      17'd18301: data = 8'h0a;
      17'd18302: data = 8'h06;
      17'd18303: data = 8'h06;
      17'd18304: data = 8'h0a;
      17'd18305: data = 8'h0a;
      17'd18306: data = 8'h0a;
      17'd18307: data = 8'h0c;
      17'd18308: data = 8'h09;
      17'd18309: data = 8'h0a;
      17'd18310: data = 8'h06;
      17'd18311: data = 8'h02;
      17'd18312: data = 8'h04;
      17'd18313: data = 8'h05;
      17'd18314: data = 8'h02;
      17'd18315: data = 8'h04;
      17'd18316: data = 8'h06;
      17'd18317: data = 8'h0c;
      17'd18318: data = 8'h0c;
      17'd18319: data = 8'h09;
      17'd18320: data = 8'h09;
      17'd18321: data = 8'h0d;
      17'd18322: data = 8'h0a;
      17'd18323: data = 8'h05;
      17'd18324: data = 8'h06;
      17'd18325: data = 8'h06;
      17'd18326: data = 8'h0a;
      17'd18327: data = 8'h0e;
      17'd18328: data = 8'h0c;
      17'd18329: data = 8'h0a;
      17'd18330: data = 8'h09;
      17'd18331: data = 8'h0a;
      17'd18332: data = 8'h0a;
      17'd18333: data = 8'h09;
      17'd18334: data = 8'h09;
      17'd18335: data = 8'h0a;
      17'd18336: data = 8'h11;
      17'd18337: data = 8'h0d;
      17'd18338: data = 8'h06;
      17'd18339: data = 8'h09;
      17'd18340: data = 8'h09;
      17'd18341: data = 8'h06;
      17'd18342: data = 8'h06;
      17'd18343: data = 8'h02;
      17'd18344: data = 8'h02;
      17'd18345: data = 8'h04;
      17'd18346: data = 8'h06;
      17'd18347: data = 8'h0a;
      17'd18348: data = 8'h05;
      17'd18349: data = 8'h04;
      17'd18350: data = 8'h05;
      17'd18351: data = 8'h02;
      17'd18352: data = 8'h00;
      17'd18353: data = 8'hfd;
      17'd18354: data = 8'hfc;
      17'd18355: data = 8'hfd;
      17'd18356: data = 8'hfd;
      17'd18357: data = 8'hfa;
      17'd18358: data = 8'hf6;
      17'd18359: data = 8'hfa;
      17'd18360: data = 8'hf9;
      17'd18361: data = 8'hf6;
      17'd18362: data = 8'hf6;
      17'd18363: data = 8'hf6;
      17'd18364: data = 8'hf9;
      17'd18365: data = 8'hf4;
      17'd18366: data = 8'hf5;
      17'd18367: data = 8'hf9;
      17'd18368: data = 8'hf5;
      17'd18369: data = 8'hf2;
      17'd18370: data = 8'hf4;
      17'd18371: data = 8'hf2;
      17'd18372: data = 8'hf1;
      17'd18373: data = 8'hf4;
      17'd18374: data = 8'hf2;
      17'd18375: data = 8'hf2;
      17'd18376: data = 8'hf5;
      17'd18377: data = 8'hf5;
      17'd18378: data = 8'hf4;
      17'd18379: data = 8'hf4;
      17'd18380: data = 8'hf6;
      17'd18381: data = 8'hf6;
      17'd18382: data = 8'hf4;
      17'd18383: data = 8'hf5;
      17'd18384: data = 8'hf9;
      17'd18385: data = 8'hf6;
      17'd18386: data = 8'hf6;
      17'd18387: data = 8'hf9;
      17'd18388: data = 8'hf9;
      17'd18389: data = 8'hf9;
      17'd18390: data = 8'hfc;
      17'd18391: data = 8'hfa;
      17'd18392: data = 8'hf9;
      17'd18393: data = 8'hfc;
      17'd18394: data = 8'hfc;
      17'd18395: data = 8'hfd;
      17'd18396: data = 8'hf6;
      17'd18397: data = 8'hfa;
      17'd18398: data = 8'h00;
      17'd18399: data = 8'hfc;
      17'd18400: data = 8'hfa;
      17'd18401: data = 8'hfd;
      17'd18402: data = 8'hfe;
      17'd18403: data = 8'hf9;
      17'd18404: data = 8'hf9;
      17'd18405: data = 8'hfa;
      17'd18406: data = 8'hfc;
      17'd18407: data = 8'hfc;
      17'd18408: data = 8'hfa;
      17'd18409: data = 8'hfa;
      17'd18410: data = 8'hfd;
      17'd18411: data = 8'hfd;
      17'd18412: data = 8'hfc;
      17'd18413: data = 8'hfc;
      17'd18414: data = 8'hfa;
      17'd18415: data = 8'hfa;
      17'd18416: data = 8'hfd;
      17'd18417: data = 8'hfa;
      17'd18418: data = 8'hfa;
      17'd18419: data = 8'hf9;
      17'd18420: data = 8'hf9;
      17'd18421: data = 8'hfc;
      17'd18422: data = 8'hfc;
      17'd18423: data = 8'hf6;
      17'd18424: data = 8'hf2;
      17'd18425: data = 8'hf9;
      17'd18426: data = 8'hfd;
      17'd18427: data = 8'hf6;
      17'd18428: data = 8'hf2;
      17'd18429: data = 8'hf4;
      17'd18430: data = 8'hf9;
      17'd18431: data = 8'hfc;
      17'd18432: data = 8'hf6;
      17'd18433: data = 8'hf5;
      17'd18434: data = 8'hf2;
      17'd18435: data = 8'hf9;
      17'd18436: data = 8'hfd;
      17'd18437: data = 8'hf6;
      17'd18438: data = 8'hf4;
      17'd18439: data = 8'hf4;
      17'd18440: data = 8'hfc;
      17'd18441: data = 8'hfa;
      17'd18442: data = 8'hf5;
      17'd18443: data = 8'hf1;
      17'd18444: data = 8'hf1;
      17'd18445: data = 8'hf2;
      17'd18446: data = 8'hf4;
      17'd18447: data = 8'hf5;
      17'd18448: data = 8'hf5;
      17'd18449: data = 8'hf2;
      17'd18450: data = 8'hef;
      17'd18451: data = 8'hf4;
      17'd18452: data = 8'hf4;
      17'd18453: data = 8'hf1;
      17'd18454: data = 8'hf4;
      17'd18455: data = 8'hf1;
      17'd18456: data = 8'hf1;
      17'd18457: data = 8'hf1;
      17'd18458: data = 8'hf1;
      17'd18459: data = 8'hf1;
      17'd18460: data = 8'hf1;
      17'd18461: data = 8'hf2;
      17'd18462: data = 8'hf4;
      17'd18463: data = 8'hf2;
      17'd18464: data = 8'hef;
      17'd18465: data = 8'hef;
      17'd18466: data = 8'hf1;
      17'd18467: data = 8'hf4;
      17'd18468: data = 8'hf5;
      17'd18469: data = 8'hf5;
      17'd18470: data = 8'hf2;
      17'd18471: data = 8'hf5;
      17'd18472: data = 8'hf9;
      17'd18473: data = 8'hf4;
      17'd18474: data = 8'hf5;
      17'd18475: data = 8'hf9;
      17'd18476: data = 8'hf5;
      17'd18477: data = 8'hf9;
      17'd18478: data = 8'hfc;
      17'd18479: data = 8'hfc;
      17'd18480: data = 8'hfa;
      17'd18481: data = 8'hf9;
      17'd18482: data = 8'hfd;
      17'd18483: data = 8'hfc;
      17'd18484: data = 8'h00;
      17'd18485: data = 8'h04;
      17'd18486: data = 8'h01;
      17'd18487: data = 8'h02;
      17'd18488: data = 8'h05;
      17'd18489: data = 8'h04;
      17'd18490: data = 8'h01;
      17'd18491: data = 8'h05;
      17'd18492: data = 8'h0c;
      17'd18493: data = 8'h06;
      17'd18494: data = 8'h0a;
      17'd18495: data = 8'h09;
      17'd18496: data = 8'h06;
      17'd18497: data = 8'h0a;
      17'd18498: data = 8'h0a;
      17'd18499: data = 8'h0c;
      17'd18500: data = 8'h09;
      17'd18501: data = 8'h0a;
      17'd18502: data = 8'h11;
      17'd18503: data = 8'h0e;
      17'd18504: data = 8'h0a;
      17'd18505: data = 8'h0e;
      17'd18506: data = 8'h12;
      17'd18507: data = 8'h11;
      17'd18508: data = 8'h0e;
      17'd18509: data = 8'h0d;
      17'd18510: data = 8'h0e;
      17'd18511: data = 8'h15;
      17'd18512: data = 8'h12;
      17'd18513: data = 8'h11;
      17'd18514: data = 8'h0d;
      17'd18515: data = 8'h0d;
      17'd18516: data = 8'h12;
      17'd18517: data = 8'h13;
      17'd18518: data = 8'h0e;
      17'd18519: data = 8'h0a;
      17'd18520: data = 8'h0d;
      17'd18521: data = 8'h0c;
      17'd18522: data = 8'h0e;
      17'd18523: data = 8'h0c;
      17'd18524: data = 8'h09;
      17'd18525: data = 8'h0a;
      17'd18526: data = 8'h0c;
      17'd18527: data = 8'h0a;
      17'd18528: data = 8'h09;
      17'd18529: data = 8'h09;
      17'd18530: data = 8'h0c;
      17'd18531: data = 8'h0c;
      17'd18532: data = 8'h09;
      17'd18533: data = 8'h09;
      17'd18534: data = 8'h0d;
      17'd18535: data = 8'h0a;
      17'd18536: data = 8'h06;
      17'd18537: data = 8'h06;
      17'd18538: data = 8'h06;
      17'd18539: data = 8'h0c;
      17'd18540: data = 8'h0a;
      17'd18541: data = 8'h05;
      17'd18542: data = 8'h06;
      17'd18543: data = 8'h0c;
      17'd18544: data = 8'h0a;
      17'd18545: data = 8'h04;
      17'd18546: data = 8'h02;
      17'd18547: data = 8'h01;
      17'd18548: data = 8'h01;
      17'd18549: data = 8'h04;
      17'd18550: data = 8'h06;
      17'd18551: data = 8'h05;
      17'd18552: data = 8'h0c;
      17'd18553: data = 8'h0d;
      17'd18554: data = 8'h06;
      17'd18555: data = 8'h06;
      17'd18556: data = 8'h0c;
      17'd18557: data = 8'h0c;
      17'd18558: data = 8'h06;
      17'd18559: data = 8'h04;
      17'd18560: data = 8'h0a;
      17'd18561: data = 8'h0c;
      17'd18562: data = 8'h0c;
      17'd18563: data = 8'h0d;
      17'd18564: data = 8'h0d;
      17'd18565: data = 8'h0a;
      17'd18566: data = 8'h0a;
      17'd18567: data = 8'h0c;
      17'd18568: data = 8'h09;
      17'd18569: data = 8'h09;
      17'd18570: data = 8'h0a;
      17'd18571: data = 8'h0d;
      17'd18572: data = 8'h0c;
      17'd18573: data = 8'h09;
      17'd18574: data = 8'h05;
      17'd18575: data = 8'h0a;
      17'd18576: data = 8'h11;
      17'd18577: data = 8'h0c;
      17'd18578: data = 8'h05;
      17'd18579: data = 8'h09;
      17'd18580: data = 8'h0a;
      17'd18581: data = 8'h0a;
      17'd18582: data = 8'h0a;
      17'd18583: data = 8'h06;
      17'd18584: data = 8'h06;
      17'd18585: data = 8'h06;
      17'd18586: data = 8'h05;
      17'd18587: data = 8'h02;
      17'd18588: data = 8'hfe;
      17'd18589: data = 8'hfe;
      17'd18590: data = 8'hfe;
      17'd18591: data = 8'hfe;
      17'd18592: data = 8'hfe;
      17'd18593: data = 8'hfd;
      17'd18594: data = 8'hfd;
      17'd18595: data = 8'hfe;
      17'd18596: data = 8'hfc;
      17'd18597: data = 8'hfa;
      17'd18598: data = 8'hf6;
      17'd18599: data = 8'hf6;
      17'd18600: data = 8'hf5;
      17'd18601: data = 8'hf6;
      17'd18602: data = 8'hf9;
      17'd18603: data = 8'hf9;
      17'd18604: data = 8'hfa;
      17'd18605: data = 8'hf9;
      17'd18606: data = 8'hf9;
      17'd18607: data = 8'hf5;
      17'd18608: data = 8'hf6;
      17'd18609: data = 8'hf6;
      17'd18610: data = 8'hf5;
      17'd18611: data = 8'hf6;
      17'd18612: data = 8'hf6;
      17'd18613: data = 8'hf4;
      17'd18614: data = 8'hf5;
      17'd18615: data = 8'hf6;
      17'd18616: data = 8'hf5;
      17'd18617: data = 8'hf5;
      17'd18618: data = 8'hf6;
      17'd18619: data = 8'hf5;
      17'd18620: data = 8'hf5;
      17'd18621: data = 8'hf9;
      17'd18622: data = 8'hfa;
      17'd18623: data = 8'hf9;
      17'd18624: data = 8'hf9;
      17'd18625: data = 8'hf9;
      17'd18626: data = 8'hf6;
      17'd18627: data = 8'hf5;
      17'd18628: data = 8'hf5;
      17'd18629: data = 8'hf6;
      17'd18630: data = 8'hfc;
      17'd18631: data = 8'hfc;
      17'd18632: data = 8'hf9;
      17'd18633: data = 8'hfc;
      17'd18634: data = 8'hfc;
      17'd18635: data = 8'hfd;
      17'd18636: data = 8'hfa;
      17'd18637: data = 8'hf5;
      17'd18638: data = 8'hf6;
      17'd18639: data = 8'hfd;
      17'd18640: data = 8'hfc;
      17'd18641: data = 8'hf9;
      17'd18642: data = 8'hfc;
      17'd18643: data = 8'hfc;
      17'd18644: data = 8'hfd;
      17'd18645: data = 8'hfc;
      17'd18646: data = 8'hfa;
      17'd18647: data = 8'hfc;
      17'd18648: data = 8'hfc;
      17'd18649: data = 8'hfd;
      17'd18650: data = 8'hfc;
      17'd18651: data = 8'hfd;
      17'd18652: data = 8'hfa;
      17'd18653: data = 8'hfa;
      17'd18654: data = 8'hfc;
      17'd18655: data = 8'hfa;
      17'd18656: data = 8'hfa;
      17'd18657: data = 8'hfa;
      17'd18658: data = 8'hfa;
      17'd18659: data = 8'hfc;
      17'd18660: data = 8'hfd;
      17'd18661: data = 8'hfd;
      17'd18662: data = 8'hfc;
      17'd18663: data = 8'hf9;
      17'd18664: data = 8'hf6;
      17'd18665: data = 8'hfc;
      17'd18666: data = 8'hfd;
      17'd18667: data = 8'hf9;
      17'd18668: data = 8'hf4;
      17'd18669: data = 8'hf6;
      17'd18670: data = 8'hf9;
      17'd18671: data = 8'hf5;
      17'd18672: data = 8'hf5;
      17'd18673: data = 8'hf5;
      17'd18674: data = 8'hf2;
      17'd18675: data = 8'hf5;
      17'd18676: data = 8'hfa;
      17'd18677: data = 8'hf4;
      17'd18678: data = 8'hf1;
      17'd18679: data = 8'hf2;
      17'd18680: data = 8'hf4;
      17'd18681: data = 8'hf6;
      17'd18682: data = 8'hf2;
      17'd18683: data = 8'hef;
      17'd18684: data = 8'hef;
      17'd18685: data = 8'hf2;
      17'd18686: data = 8'hef;
      17'd18687: data = 8'hef;
      17'd18688: data = 8'hf1;
      17'd18689: data = 8'hed;
      17'd18690: data = 8'hec;
      17'd18691: data = 8'hef;
      17'd18692: data = 8'hef;
      17'd18693: data = 8'hef;
      17'd18694: data = 8'hef;
      17'd18695: data = 8'hec;
      17'd18696: data = 8'hed;
      17'd18697: data = 8'hef;
      17'd18698: data = 8'hed;
      17'd18699: data = 8'hec;
      17'd18700: data = 8'hec;
      17'd18701: data = 8'hec;
      17'd18702: data = 8'hf1;
      17'd18703: data = 8'hf1;
      17'd18704: data = 8'hef;
      17'd18705: data = 8'hef;
      17'd18706: data = 8'hed;
      17'd18707: data = 8'hef;
      17'd18708: data = 8'hf1;
      17'd18709: data = 8'hf1;
      17'd18710: data = 8'hf2;
      17'd18711: data = 8'hf5;
      17'd18712: data = 8'hf4;
      17'd18713: data = 8'hf5;
      17'd18714: data = 8'hf5;
      17'd18715: data = 8'hf4;
      17'd18716: data = 8'hf4;
      17'd18717: data = 8'hf6;
      17'd18718: data = 8'hf6;
      17'd18719: data = 8'hf9;
      17'd18720: data = 8'hfa;
      17'd18721: data = 8'hfa;
      17'd18722: data = 8'hfc;
      17'd18723: data = 8'hfe;
      17'd18724: data = 8'hfe;
      17'd18725: data = 8'h00;
      17'd18726: data = 8'hfe;
      17'd18727: data = 8'h00;
      17'd18728: data = 8'h02;
      17'd18729: data = 8'h06;
      17'd18730: data = 8'h05;
      17'd18731: data = 8'h00;
      17'd18732: data = 8'h04;
      17'd18733: data = 8'h0c;
      17'd18734: data = 8'h0c;
      17'd18735: data = 8'h06;
      17'd18736: data = 8'h04;
      17'd18737: data = 8'h05;
      17'd18738: data = 8'h0c;
      17'd18739: data = 8'h0c;
      17'd18740: data = 8'h0a;
      17'd18741: data = 8'h05;
      17'd18742: data = 8'h06;
      17'd18743: data = 8'h11;
      17'd18744: data = 8'h12;
      17'd18745: data = 8'h0c;
      17'd18746: data = 8'h09;
      17'd18747: data = 8'h0d;
      17'd18748: data = 8'h12;
      17'd18749: data = 8'h15;
      17'd18750: data = 8'h0e;
      17'd18751: data = 8'h0d;
      17'd18752: data = 8'h0e;
      17'd18753: data = 8'h13;
      17'd18754: data = 8'h0e;
      17'd18755: data = 8'h0d;
      17'd18756: data = 8'h0c;
      17'd18757: data = 8'h0d;
      17'd18758: data = 8'h13;
      17'd18759: data = 8'h0e;
      17'd18760: data = 8'h0a;
      17'd18761: data = 8'h0e;
      17'd18762: data = 8'h11;
      17'd18763: data = 8'h0d;
      17'd18764: data = 8'h11;
      17'd18765: data = 8'h0c;
      17'd18766: data = 8'h0c;
      17'd18767: data = 8'h0a;
      17'd18768: data = 8'h0e;
      17'd18769: data = 8'h0a;
      17'd18770: data = 8'h0c;
      17'd18771: data = 8'h0d;
      17'd18772: data = 8'h0d;
      17'd18773: data = 8'h06;
      17'd18774: data = 8'h06;
      17'd18775: data = 8'h0c;
      17'd18776: data = 8'h09;
      17'd18777: data = 8'h09;
      17'd18778: data = 8'h09;
      17'd18779: data = 8'h0d;
      17'd18780: data = 8'h0e;
      17'd18781: data = 8'h0c;
      17'd18782: data = 8'h05;
      17'd18783: data = 8'h02;
      17'd18784: data = 8'h04;
      17'd18785: data = 8'h02;
      17'd18786: data = 8'h01;
      17'd18787: data = 8'h01;
      17'd18788: data = 8'h01;
      17'd18789: data = 8'h0a;
      17'd18790: data = 8'h0d;
      17'd18791: data = 8'h06;
      17'd18792: data = 8'h05;
      17'd18793: data = 8'h09;
      17'd18794: data = 8'h09;
      17'd18795: data = 8'h06;
      17'd18796: data = 8'h09;
      17'd18797: data = 8'h05;
      17'd18798: data = 8'h06;
      17'd18799: data = 8'h06;
      17'd18800: data = 8'h0d;
      17'd18801: data = 8'h0c;
      17'd18802: data = 8'h04;
      17'd18803: data = 8'h06;
      17'd18804: data = 8'h09;
      17'd18805: data = 8'h0d;
      17'd18806: data = 8'h09;
      17'd18807: data = 8'h09;
      17'd18808: data = 8'h0d;
      17'd18809: data = 8'h0c;
      17'd18810: data = 8'h0d;
      17'd18811: data = 8'h0c;
      17'd18812: data = 8'h0a;
      17'd18813: data = 8'h09;
      17'd18814: data = 8'h06;
      17'd18815: data = 8'h04;
      17'd18816: data = 8'h05;
      17'd18817: data = 8'h0a;
      17'd18818: data = 8'h0a;
      17'd18819: data = 8'h09;
      17'd18820: data = 8'h0c;
      17'd18821: data = 8'h0c;
      17'd18822: data = 8'h09;
      17'd18823: data = 8'h09;
      17'd18824: data = 8'h06;
      17'd18825: data = 8'h02;
      17'd18826: data = 8'h01;
      17'd18827: data = 8'h04;
      17'd18828: data = 8'h00;
      17'd18829: data = 8'hfd;
      17'd18830: data = 8'hfe;
      17'd18831: data = 8'hfd;
      17'd18832: data = 8'h00;
      17'd18833: data = 8'hfe;
      17'd18834: data = 8'hf9;
      17'd18835: data = 8'hfa;
      17'd18836: data = 8'hfa;
      17'd18837: data = 8'hfa;
      17'd18838: data = 8'hfc;
      17'd18839: data = 8'hf9;
      17'd18840: data = 8'hf6;
      17'd18841: data = 8'hf6;
      17'd18842: data = 8'hf9;
      17'd18843: data = 8'hf6;
      17'd18844: data = 8'hf2;
      17'd18845: data = 8'hf2;
      17'd18846: data = 8'hf6;
      17'd18847: data = 8'hf6;
      17'd18848: data = 8'hf9;
      17'd18849: data = 8'hf9;
      17'd18850: data = 8'hf6;
      17'd18851: data = 8'hfa;
      17'd18852: data = 8'hfa;
      17'd18853: data = 8'hf5;
      17'd18854: data = 8'hf6;
      17'd18855: data = 8'hf4;
      17'd18856: data = 8'hf5;
      17'd18857: data = 8'hf6;
      17'd18858: data = 8'hf4;
      17'd18859: data = 8'hf9;
      17'd18860: data = 8'hfa;
      17'd18861: data = 8'hfc;
      17'd18862: data = 8'hfc;
      17'd18863: data = 8'hfc;
      17'd18864: data = 8'hfc;
      17'd18865: data = 8'hfd;
      17'd18866: data = 8'hfd;
      17'd18867: data = 8'hfa;
      17'd18868: data = 8'hfa;
      17'd18869: data = 8'hfd;
      17'd18870: data = 8'h01;
      17'd18871: data = 8'h00;
      17'd18872: data = 8'hfc;
      17'd18873: data = 8'hfc;
      17'd18874: data = 8'hfc;
      17'd18875: data = 8'hfe;
      17'd18876: data = 8'h00;
      17'd18877: data = 8'hf9;
      17'd18878: data = 8'hfa;
      17'd18879: data = 8'h00;
      17'd18880: data = 8'h00;
      17'd18881: data = 8'hfd;
      17'd18882: data = 8'hfd;
      17'd18883: data = 8'hfe;
      17'd18884: data = 8'hfe;
      17'd18885: data = 8'hfc;
      17'd18886: data = 8'hf6;
      17'd18887: data = 8'hf9;
      17'd18888: data = 8'hfc;
      17'd18889: data = 8'hfd;
      17'd18890: data = 8'hfd;
      17'd18891: data = 8'hfc;
      17'd18892: data = 8'hfd;
      17'd18893: data = 8'hfd;
      17'd18894: data = 8'hfc;
      17'd18895: data = 8'hfc;
      17'd18896: data = 8'hfa;
      17'd18897: data = 8'hf6;
      17'd18898: data = 8'hfa;
      17'd18899: data = 8'hfa;
      17'd18900: data = 8'hf6;
      17'd18901: data = 8'hf9;
      17'd18902: data = 8'hfc;
      17'd18903: data = 8'hfc;
      17'd18904: data = 8'hfa;
      17'd18905: data = 8'hf9;
      17'd18906: data = 8'hf6;
      17'd18907: data = 8'hf5;
      17'd18908: data = 8'hfa;
      17'd18909: data = 8'hf6;
      17'd18910: data = 8'hf5;
      17'd18911: data = 8'hf9;
      17'd18912: data = 8'hfa;
      17'd18913: data = 8'hf4;
      17'd18914: data = 8'hf1;
      17'd18915: data = 8'hf1;
      17'd18916: data = 8'hf2;
      17'd18917: data = 8'hf4;
      17'd18918: data = 8'hf2;
      17'd18919: data = 8'hf1;
      17'd18920: data = 8'hf4;
      17'd18921: data = 8'hf4;
      17'd18922: data = 8'hf4;
      17'd18923: data = 8'hf2;
      17'd18924: data = 8'hef;
      17'd18925: data = 8'hec;
      17'd18926: data = 8'hed;
      17'd18927: data = 8'hed;
      17'd18928: data = 8'hed;
      17'd18929: data = 8'hf2;
      17'd18930: data = 8'hf1;
      17'd18931: data = 8'hed;
      17'd18932: data = 8'hed;
      17'd18933: data = 8'hf2;
      17'd18934: data = 8'hf1;
      17'd18935: data = 8'hed;
      17'd18936: data = 8'hed;
      17'd18937: data = 8'hf1;
      17'd18938: data = 8'hf2;
      17'd18939: data = 8'hf1;
      17'd18940: data = 8'hef;
      17'd18941: data = 8'hf1;
      17'd18942: data = 8'hef;
      17'd18943: data = 8'hef;
      17'd18944: data = 8'hf2;
      17'd18945: data = 8'hf2;
      17'd18946: data = 8'hf2;
      17'd18947: data = 8'hf5;
      17'd18948: data = 8'hf4;
      17'd18949: data = 8'hf2;
      17'd18950: data = 8'hf4;
      17'd18951: data = 8'hf9;
      17'd18952: data = 8'hf9;
      17'd18953: data = 8'hf4;
      17'd18954: data = 8'hf5;
      17'd18955: data = 8'hf9;
      17'd18956: data = 8'hfa;
      17'd18957: data = 8'hfa;
      17'd18958: data = 8'hfa;
      17'd18959: data = 8'hfc;
      17'd18960: data = 8'hfc;
      17'd18961: data = 8'hfe;
      17'd18962: data = 8'h01;
      17'd18963: data = 8'h02;
      17'd18964: data = 8'h01;
      17'd18965: data = 8'h02;
      17'd18966: data = 8'h05;
      17'd18967: data = 8'h01;
      17'd18968: data = 8'h02;
      17'd18969: data = 8'h06;
      17'd18970: data = 8'h04;
      17'd18971: data = 8'h05;
      17'd18972: data = 8'h09;
      17'd18973: data = 8'h09;
      17'd18974: data = 8'h0a;
      17'd18975: data = 8'h0c;
      17'd18976: data = 8'h0d;
      17'd18977: data = 8'h0c;
      17'd18978: data = 8'h0c;
      17'd18979: data = 8'h0e;
      17'd18980: data = 8'h0d;
      17'd18981: data = 8'h0d;
      17'd18982: data = 8'h11;
      17'd18983: data = 8'h0e;
      17'd18984: data = 8'h0e;
      17'd18985: data = 8'h0d;
      17'd18986: data = 8'h0e;
      17'd18987: data = 8'h12;
      17'd18988: data = 8'h13;
      17'd18989: data = 8'h11;
      17'd18990: data = 8'h0e;
      17'd18991: data = 8'h13;
      17'd18992: data = 8'h13;
      17'd18993: data = 8'h12;
      17'd18994: data = 8'h12;
      17'd18995: data = 8'h0e;
      17'd18996: data = 8'h0e;
      17'd18997: data = 8'h11;
      17'd18998: data = 8'h12;
      17'd18999: data = 8'h0e;
      17'd19000: data = 8'h0d;
      17'd19001: data = 8'h0e;
      17'd19002: data = 8'h0e;
      17'd19003: data = 8'h11;
      17'd19004: data = 8'h11;
      17'd19005: data = 8'h0d;
      17'd19006: data = 8'h0d;
      17'd19007: data = 8'h0e;
      17'd19008: data = 8'h0c;
      17'd19009: data = 8'h0a;
      17'd19010: data = 8'h0a;
      17'd19011: data = 8'h0a;
      17'd19012: data = 8'h09;
      17'd19013: data = 8'h06;
      17'd19014: data = 8'h09;
      17'd19015: data = 8'h09;
      17'd19016: data = 8'h09;
      17'd19017: data = 8'h0a;
      17'd19018: data = 8'h0a;
      17'd19019: data = 8'h09;
      17'd19020: data = 8'h04;
      17'd19021: data = 8'h02;
      17'd19022: data = 8'h02;
      17'd19023: data = 8'h00;
      17'd19024: data = 8'h00;
      17'd19025: data = 8'h02;
      17'd19026: data = 8'h06;
      17'd19027: data = 8'h04;
      17'd19028: data = 8'h02;
      17'd19029: data = 8'h04;
      17'd19030: data = 8'h02;
      17'd19031: data = 8'h04;
      17'd19032: data = 8'h05;
      17'd19033: data = 8'h04;
      17'd19034: data = 8'h05;
      17'd19035: data = 8'h06;
      17'd19036: data = 8'h05;
      17'd19037: data = 8'h05;
      17'd19038: data = 8'h09;
      17'd19039: data = 8'h06;
      17'd19040: data = 8'h04;
      17'd19041: data = 8'h05;
      17'd19042: data = 8'h04;
      17'd19043: data = 8'h05;
      17'd19044: data = 8'h06;
      17'd19045: data = 8'h04;
      17'd19046: data = 8'h09;
      17'd19047: data = 8'h0c;
      17'd19048: data = 8'h0a;
      17'd19049: data = 8'h0d;
      17'd19050: data = 8'h0d;
      17'd19051: data = 8'h06;
      17'd19052: data = 8'h09;
      17'd19053: data = 8'h0c;
      17'd19054: data = 8'h09;
      17'd19055: data = 8'h05;
      17'd19056: data = 8'h06;
      17'd19057: data = 8'h09;
      17'd19058: data = 8'h0a;
      17'd19059: data = 8'h0d;
      17'd19060: data = 8'h09;
      17'd19061: data = 8'h05;
      17'd19062: data = 8'h06;
      17'd19063: data = 8'h02;
      17'd19064: data = 8'h04;
      17'd19065: data = 8'h01;
      17'd19066: data = 8'hfd;
      17'd19067: data = 8'h00;
      17'd19068: data = 8'h01;
      17'd19069: data = 8'hfe;
      17'd19070: data = 8'hfa;
      17'd19071: data = 8'hf9;
      17'd19072: data = 8'hfa;
      17'd19073: data = 8'hfc;
      17'd19074: data = 8'hfc;
      17'd19075: data = 8'hfa;
      17'd19076: data = 8'hfd;
      17'd19077: data = 8'hfe;
      17'd19078: data = 8'hfd;
      17'd19079: data = 8'hfc;
      17'd19080: data = 8'hfa;
      17'd19081: data = 8'hf9;
      17'd19082: data = 8'hf4;
      17'd19083: data = 8'hf2;
      17'd19084: data = 8'hf4;
      17'd19085: data = 8'hf4;
      17'd19086: data = 8'hf5;
      17'd19087: data = 8'hf9;
      17'd19088: data = 8'hf9;
      17'd19089: data = 8'hfa;
      17'd19090: data = 8'hfa;
      17'd19091: data = 8'hf6;
      17'd19092: data = 8'hfa;
      17'd19093: data = 8'hf9;
      17'd19094: data = 8'hf5;
      17'd19095: data = 8'hf4;
      17'd19096: data = 8'hf4;
      17'd19097: data = 8'hf6;
      17'd19098: data = 8'hf5;
      17'd19099: data = 8'hf5;
      17'd19100: data = 8'hf9;
      17'd19101: data = 8'hfc;
      17'd19102: data = 8'hfa;
      17'd19103: data = 8'hfa;
      17'd19104: data = 8'hfc;
      17'd19105: data = 8'hfc;
      17'd19106: data = 8'hfd;
      17'd19107: data = 8'hfc;
      17'd19108: data = 8'hfe;
      17'd19109: data = 8'hfe;
      17'd19110: data = 8'hfc;
      17'd19111: data = 8'hfa;
      17'd19112: data = 8'hf6;
      17'd19113: data = 8'hf6;
      17'd19114: data = 8'hf6;
      17'd19115: data = 8'hfa;
      17'd19116: data = 8'hfa;
      17'd19117: data = 8'hfc;
      17'd19118: data = 8'h01;
      17'd19119: data = 8'h02;
      17'd19120: data = 8'h00;
      17'd19121: data = 8'hfe;
      17'd19122: data = 8'hfe;
      17'd19123: data = 8'hfd;
      17'd19124: data = 8'hfc;
      17'd19125: data = 8'hfc;
      17'd19126: data = 8'hfc;
      17'd19127: data = 8'hfd;
      17'd19128: data = 8'hfc;
      17'd19129: data = 8'hfc;
      17'd19130: data = 8'hfe;
      17'd19131: data = 8'hfd;
      17'd19132: data = 8'hfd;
      17'd19133: data = 8'hfd;
      17'd19134: data = 8'hfd;
      17'd19135: data = 8'hfd;
      17'd19136: data = 8'hfd;
      17'd19137: data = 8'hfc;
      17'd19138: data = 8'hfa;
      17'd19139: data = 8'hfa;
      17'd19140: data = 8'hfa;
      17'd19141: data = 8'hf6;
      17'd19142: data = 8'hfa;
      17'd19143: data = 8'hf9;
      17'd19144: data = 8'hf4;
      17'd19145: data = 8'hf6;
      17'd19146: data = 8'hf6;
      17'd19147: data = 8'hf9;
      17'd19148: data = 8'hf9;
      17'd19149: data = 8'hf6;
      17'd19150: data = 8'hf9;
      17'd19151: data = 8'hfc;
      17'd19152: data = 8'hf6;
      17'd19153: data = 8'hf2;
      17'd19154: data = 8'hef;
      17'd19155: data = 8'hef;
      17'd19156: data = 8'hef;
      17'd19157: data = 8'hef;
      17'd19158: data = 8'hed;
      17'd19159: data = 8'hed;
      17'd19160: data = 8'hef;
      17'd19161: data = 8'hed;
      17'd19162: data = 8'hf1;
      17'd19163: data = 8'hec;
      17'd19164: data = 8'heb;
      17'd19165: data = 8'hec;
      17'd19166: data = 8'hec;
      17'd19167: data = 8'hec;
      17'd19168: data = 8'hec;
      17'd19169: data = 8'hec;
      17'd19170: data = 8'hec;
      17'd19171: data = 8'he9;
      17'd19172: data = 8'he9;
      17'd19173: data = 8'heb;
      17'd19174: data = 8'heb;
      17'd19175: data = 8'heb;
      17'd19176: data = 8'hec;
      17'd19177: data = 8'heb;
      17'd19178: data = 8'hed;
      17'd19179: data = 8'hf2;
      17'd19180: data = 8'hef;
      17'd19181: data = 8'hec;
      17'd19182: data = 8'hef;
      17'd19183: data = 8'hed;
      17'd19184: data = 8'hed;
      17'd19185: data = 8'hf1;
      17'd19186: data = 8'hef;
      17'd19187: data = 8'hf1;
      17'd19188: data = 8'hf2;
      17'd19189: data = 8'hf4;
      17'd19190: data = 8'hf6;
      17'd19191: data = 8'hf5;
      17'd19192: data = 8'hf6;
      17'd19193: data = 8'hf6;
      17'd19194: data = 8'hfa;
      17'd19195: data = 8'hf9;
      17'd19196: data = 8'hfa;
      17'd19197: data = 8'hfc;
      17'd19198: data = 8'hfa;
      17'd19199: data = 8'hfc;
      17'd19200: data = 8'hfd;
      17'd19201: data = 8'h02;
      17'd19202: data = 8'h02;
      17'd19203: data = 8'h01;
      17'd19204: data = 8'h04;
      17'd19205: data = 8'h06;
      17'd19206: data = 8'h04;
      17'd19207: data = 8'h02;
      17'd19208: data = 8'h09;
      17'd19209: data = 8'h0a;
      17'd19210: data = 8'h06;
      17'd19211: data = 8'h0c;
      17'd19212: data = 8'h0e;
      17'd19213: data = 8'h11;
      17'd19214: data = 8'h0e;
      17'd19215: data = 8'h0d;
      17'd19216: data = 8'h0e;
      17'd19217: data = 8'h11;
      17'd19218: data = 8'h15;
      17'd19219: data = 8'h13;
      17'd19220: data = 8'h12;
      17'd19221: data = 8'h15;
      17'd19222: data = 8'h16;
      17'd19223: data = 8'h16;
      17'd19224: data = 8'h16;
      17'd19225: data = 8'h15;
      17'd19226: data = 8'h15;
      17'd19227: data = 8'h19;
      17'd19228: data = 8'h19;
      17'd19229: data = 8'h13;
      17'd19230: data = 8'h15;
      17'd19231: data = 8'h19;
      17'd19232: data = 8'h15;
      17'd19233: data = 8'h13;
      17'd19234: data = 8'h13;
      17'd19235: data = 8'h16;
      17'd19236: data = 8'h15;
      17'd19237: data = 8'h13;
      17'd19238: data = 8'h15;
      17'd19239: data = 8'h12;
      17'd19240: data = 8'h15;
      17'd19241: data = 8'h13;
      17'd19242: data = 8'h12;
      17'd19243: data = 8'h11;
      17'd19244: data = 8'h0e;
      17'd19245: data = 8'h11;
      17'd19246: data = 8'h0c;
      17'd19247: data = 8'h0a;
      17'd19248: data = 8'h09;
      17'd19249: data = 8'h0a;
      17'd19250: data = 8'h0a;
      17'd19251: data = 8'h09;
      17'd19252: data = 8'h06;
      17'd19253: data = 8'h05;
      17'd19254: data = 8'h05;
      17'd19255: data = 8'h09;
      17'd19256: data = 8'h02;
      17'd19257: data = 8'hfd;
      17'd19258: data = 8'h00;
      17'd19259: data = 8'h01;
      17'd19260: data = 8'h02;
      17'd19261: data = 8'hfe;
      17'd19262: data = 8'hfe;
      17'd19263: data = 8'h02;
      17'd19264: data = 8'h04;
      17'd19265: data = 8'h01;
      17'd19266: data = 8'hfe;
      17'd19267: data = 8'hfe;
      17'd19268: data = 8'h01;
      17'd19269: data = 8'h02;
      17'd19270: data = 8'h04;
      17'd19271: data = 8'h02;
      17'd19272: data = 8'h01;
      17'd19273: data = 8'h05;
      17'd19274: data = 8'h06;
      17'd19275: data = 8'h06;
      17'd19276: data = 8'h01;
      17'd19277: data = 8'h01;
      17'd19278: data = 8'h05;
      17'd19279: data = 8'h05;
      17'd19280: data = 8'h06;
      17'd19281: data = 8'h06;
      17'd19282: data = 8'h06;
      17'd19283: data = 8'h0a;
      17'd19284: data = 8'h0a;
      17'd19285: data = 8'h09;
      17'd19286: data = 8'h0a;
      17'd19287: data = 8'h0d;
      17'd19288: data = 8'h0c;
      17'd19289: data = 8'h0a;
      17'd19290: data = 8'h0a;
      17'd19291: data = 8'h0a;
      17'd19292: data = 8'h0a;
      17'd19293: data = 8'h0a;
      17'd19294: data = 8'h0d;
      17'd19295: data = 8'h0c;
      17'd19296: data = 8'h0a;
      17'd19297: data = 8'h06;
      17'd19298: data = 8'h05;
      17'd19299: data = 8'h06;
      17'd19300: data = 8'h04;
      17'd19301: data = 8'h02;
      17'd19302: data = 8'h02;
      17'd19303: data = 8'h01;
      17'd19304: data = 8'h00;
      17'd19305: data = 8'hfd;
      17'd19306: data = 8'hfd;
      17'd19307: data = 8'hfa;
      17'd19308: data = 8'hf9;
      17'd19309: data = 8'hfc;
      17'd19310: data = 8'hf9;
      17'd19311: data = 8'hf9;
      17'd19312: data = 8'hfc;
      17'd19313: data = 8'hfa;
      17'd19314: data = 8'hf9;
      17'd19315: data = 8'hfc;
      17'd19316: data = 8'hfa;
      17'd19317: data = 8'hfa;
      17'd19318: data = 8'hf9;
      17'd19319: data = 8'hf2;
      17'd19320: data = 8'hf2;
      17'd19321: data = 8'hf4;
      17'd19322: data = 8'hf2;
      17'd19323: data = 8'hf4;
      17'd19324: data = 8'hf6;
      17'd19325: data = 8'hf9;
      17'd19326: data = 8'hf6;
      17'd19327: data = 8'hf5;
      17'd19328: data = 8'hf9;
      17'd19329: data = 8'hf6;
      17'd19330: data = 8'hf5;
      17'd19331: data = 8'hf9;
      17'd19332: data = 8'hf9;
      17'd19333: data = 8'hfa;
      17'd19334: data = 8'hfe;
      17'd19335: data = 8'hfd;
      17'd19336: data = 8'hfc;
      17'd19337: data = 8'hfc;
      17'd19338: data = 8'hfc;
      17'd19339: data = 8'hfc;
      17'd19340: data = 8'hfe;
      17'd19341: data = 8'h00;
      17'd19342: data = 8'hfe;
      17'd19343: data = 8'h00;
      17'd19344: data = 8'h02;
      17'd19345: data = 8'h01;
      17'd19346: data = 8'hfe;
      17'd19347: data = 8'h01;
      17'd19348: data = 8'hfe;
      17'd19349: data = 8'hfc;
      17'd19350: data = 8'hfc;
      17'd19351: data = 8'hfc;
      17'd19352: data = 8'h00;
      17'd19353: data = 8'hfd;
      17'd19354: data = 8'hfd;
      17'd19355: data = 8'hfd;
      17'd19356: data = 8'hfd;
      17'd19357: data = 8'h01;
      17'd19358: data = 8'h01;
      17'd19359: data = 8'hfe;
      17'd19360: data = 8'h01;
      17'd19361: data = 8'h05;
      17'd19362: data = 8'h01;
      17'd19363: data = 8'hfd;
      17'd19364: data = 8'hfd;
      17'd19365: data = 8'hfd;
      17'd19366: data = 8'hfe;
      17'd19367: data = 8'hfe;
      17'd19368: data = 8'hfc;
      17'd19369: data = 8'hfa;
      17'd19370: data = 8'hfd;
      17'd19371: data = 8'hfc;
      17'd19372: data = 8'hf9;
      17'd19373: data = 8'hf9;
      17'd19374: data = 8'hf9;
      17'd19375: data = 8'hf9;
      17'd19376: data = 8'hfc;
      17'd19377: data = 8'hfd;
      17'd19378: data = 8'hf6;
      17'd19379: data = 8'hf6;
      17'd19380: data = 8'hfa;
      17'd19381: data = 8'hfa;
      17'd19382: data = 8'hf6;
      17'd19383: data = 8'hf5;
      17'd19384: data = 8'hf4;
      17'd19385: data = 8'hf6;
      17'd19386: data = 8'hfa;
      17'd19387: data = 8'hf9;
      17'd19388: data = 8'hf4;
      17'd19389: data = 8'hf4;
      17'd19390: data = 8'hf4;
      17'd19391: data = 8'hf2;
      17'd19392: data = 8'hf2;
      17'd19393: data = 8'hf1;
      17'd19394: data = 8'hf1;
      17'd19395: data = 8'hf1;
      17'd19396: data = 8'hec;
      17'd19397: data = 8'heb;
      17'd19398: data = 8'hec;
      17'd19399: data = 8'he9;
      17'd19400: data = 8'heb;
      17'd19401: data = 8'hec;
      17'd19402: data = 8'heb;
      17'd19403: data = 8'heb;
      17'd19404: data = 8'hed;
      17'd19405: data = 8'heb;
      17'd19406: data = 8'he9;
      17'd19407: data = 8'hec;
      17'd19408: data = 8'he9;
      17'd19409: data = 8'he9;
      17'd19410: data = 8'he9;
      17'd19411: data = 8'he7;
      17'd19412: data = 8'he7;
      17'd19413: data = 8'hec;
      17'd19414: data = 8'hef;
      17'd19415: data = 8'hed;
      17'd19416: data = 8'hec;
      17'd19417: data = 8'he7;
      17'd19418: data = 8'he7;
      17'd19419: data = 8'hed;
      17'd19420: data = 8'hf1;
      17'd19421: data = 8'hf2;
      17'd19422: data = 8'hef;
      17'd19423: data = 8'hed;
      17'd19424: data = 8'hec;
      17'd19425: data = 8'hec;
      17'd19426: data = 8'hed;
      17'd19427: data = 8'hf1;
      17'd19428: data = 8'hf4;
      17'd19429: data = 8'hf6;
      17'd19430: data = 8'hf6;
      17'd19431: data = 8'hf5;
      17'd19432: data = 8'hf6;
      17'd19433: data = 8'hf9;
      17'd19434: data = 8'h00;
      17'd19435: data = 8'h04;
      17'd19436: data = 8'h00;
      17'd19437: data = 8'hfd;
      17'd19438: data = 8'h00;
      17'd19439: data = 8'h02;
      17'd19440: data = 8'h06;
      17'd19441: data = 8'h05;
      17'd19442: data = 8'h04;
      17'd19443: data = 8'h05;
      17'd19444: data = 8'h0a;
      17'd19445: data = 8'h0d;
      17'd19446: data = 8'h0a;
      17'd19447: data = 8'h0c;
      17'd19448: data = 8'h0c;
      17'd19449: data = 8'h12;
      17'd19450: data = 8'h11;
      17'd19451: data = 8'h0d;
      17'd19452: data = 8'h0e;
      17'd19453: data = 8'h13;
      17'd19454: data = 8'h15;
      17'd19455: data = 8'h13;
      17'd19456: data = 8'h15;
      17'd19457: data = 8'h16;
      17'd19458: data = 8'h13;
      17'd19459: data = 8'h11;
      17'd19460: data = 8'h15;
      17'd19461: data = 8'h1a;
      17'd19462: data = 8'h1a;
      17'd19463: data = 8'h19;
      17'd19464: data = 8'h16;
      17'd19465: data = 8'h13;
      17'd19466: data = 8'h19;
      17'd19467: data = 8'h15;
      17'd19468: data = 8'h15;
      17'd19469: data = 8'h16;
      17'd19470: data = 8'h15;
      17'd19471: data = 8'h15;
      17'd19472: data = 8'h15;
      17'd19473: data = 8'h15;
      17'd19474: data = 8'h11;
      17'd19475: data = 8'h12;
      17'd19476: data = 8'h11;
      17'd19477: data = 8'h11;
      17'd19478: data = 8'h12;
      17'd19479: data = 8'h11;
      17'd19480: data = 8'h0e;
      17'd19481: data = 8'h0e;
      17'd19482: data = 8'h0e;
      17'd19483: data = 8'h0a;
      17'd19484: data = 8'h06;
      17'd19485: data = 8'h0c;
      17'd19486: data = 8'h0a;
      17'd19487: data = 8'h05;
      17'd19488: data = 8'h04;
      17'd19489: data = 8'h04;
      17'd19490: data = 8'h04;
      17'd19491: data = 8'h01;
      17'd19492: data = 8'h00;
      17'd19493: data = 8'h01;
      17'd19494: data = 8'h02;
      17'd19495: data = 8'h01;
      17'd19496: data = 8'h00;
      17'd19497: data = 8'h01;
      17'd19498: data = 8'h02;
      17'd19499: data = 8'h02;
      17'd19500: data = 8'hfe;
      17'd19501: data = 8'hfd;
      17'd19502: data = 8'h01;
      17'd19503: data = 8'h02;
      17'd19504: data = 8'h00;
      17'd19505: data = 8'h04;
      17'd19506: data = 8'h06;
      17'd19507: data = 8'h05;
      17'd19508: data = 8'h05;
      17'd19509: data = 8'h05;
      17'd19510: data = 8'h05;
      17'd19511: data = 8'h05;
      17'd19512: data = 8'h05;
      17'd19513: data = 8'h06;
      17'd19514: data = 8'h06;
      17'd19515: data = 8'h06;
      17'd19516: data = 8'h06;
      17'd19517: data = 8'h0d;
      17'd19518: data = 8'h0d;
      17'd19519: data = 8'h0a;
      17'd19520: data = 8'h0a;
      17'd19521: data = 8'h0d;
      17'd19522: data = 8'h0e;
      17'd19523: data = 8'h0e;
      17'd19524: data = 8'h0d;
      17'd19525: data = 8'h0c;
      17'd19526: data = 8'h0d;
      17'd19527: data = 8'h0e;
      17'd19528: data = 8'h0a;
      17'd19529: data = 8'h0a;
      17'd19530: data = 8'h0a;
      17'd19531: data = 8'h06;
      17'd19532: data = 8'h04;
      17'd19533: data = 8'h01;
      17'd19534: data = 8'h00;
      17'd19535: data = 8'h02;
      17'd19536: data = 8'h00;
      17'd19537: data = 8'h00;
      17'd19538: data = 8'h00;
      17'd19539: data = 8'hfe;
      17'd19540: data = 8'hfc;
      17'd19541: data = 8'hf9;
      17'd19542: data = 8'hf9;
      17'd19543: data = 8'hf5;
      17'd19544: data = 8'hf5;
      17'd19545: data = 8'hf4;
      17'd19546: data = 8'hf6;
      17'd19547: data = 8'hf5;
      17'd19548: data = 8'hf6;
      17'd19549: data = 8'hf6;
      17'd19550: data = 8'hf5;
      17'd19551: data = 8'hf5;
      17'd19552: data = 8'hf6;
      17'd19553: data = 8'hf5;
      17'd19554: data = 8'hf2;
      17'd19555: data = 8'hf2;
      17'd19556: data = 8'hf4;
      17'd19557: data = 8'hf4;
      17'd19558: data = 8'hf2;
      17'd19559: data = 8'hf6;
      17'd19560: data = 8'hf6;
      17'd19561: data = 8'hf4;
      17'd19562: data = 8'hf4;
      17'd19563: data = 8'hf9;
      17'd19564: data = 8'hf9;
      17'd19565: data = 8'hf9;
      17'd19566: data = 8'hfa;
      17'd19567: data = 8'hfc;
      17'd19568: data = 8'hfd;
      17'd19569: data = 8'hfe;
      17'd19570: data = 8'h01;
      17'd19571: data = 8'hfe;
      17'd19572: data = 8'hfd;
      17'd19573: data = 8'h01;
      17'd19574: data = 8'h01;
      17'd19575: data = 8'h00;
      17'd19576: data = 8'h01;
      17'd19577: data = 8'h02;
      17'd19578: data = 8'h02;
      17'd19579: data = 8'h02;
      17'd19580: data = 8'h06;
      17'd19581: data = 8'h05;
      17'd19582: data = 8'h02;
      17'd19583: data = 8'h02;
      17'd19584: data = 8'h02;
      17'd19585: data = 8'h02;
      17'd19586: data = 8'h00;
      17'd19587: data = 8'h00;
      17'd19588: data = 8'hfe;
      17'd19589: data = 8'h01;
      17'd19590: data = 8'h01;
      17'd19591: data = 8'h00;
      17'd19592: data = 8'h02;
      17'd19593: data = 8'h01;
      17'd19594: data = 8'h00;
      17'd19595: data = 8'h00;
      17'd19596: data = 8'h00;
      17'd19597: data = 8'hfe;
      17'd19598: data = 8'hfe;
      17'd19599: data = 8'h01;
      17'd19600: data = 8'hfd;
      17'd19601: data = 8'hfd;
      17'd19602: data = 8'hfe;
      17'd19603: data = 8'hfa;
      17'd19604: data = 8'hfa;
      17'd19605: data = 8'hfc;
      17'd19606: data = 8'hf9;
      17'd19607: data = 8'hf4;
      17'd19608: data = 8'hf6;
      17'd19609: data = 8'hfa;
      17'd19610: data = 8'hf9;
      17'd19611: data = 8'hfa;
      17'd19612: data = 8'hf6;
      17'd19613: data = 8'hf4;
      17'd19614: data = 8'hf4;
      17'd19615: data = 8'hf5;
      17'd19616: data = 8'hf6;
      17'd19617: data = 8'hf5;
      17'd19618: data = 8'hf4;
      17'd19619: data = 8'hf4;
      17'd19620: data = 8'hf6;
      17'd19621: data = 8'hf5;
      17'd19622: data = 8'hf2;
      17'd19623: data = 8'hf4;
      17'd19624: data = 8'hf4;
      17'd19625: data = 8'hf1;
      17'd19626: data = 8'hed;
      17'd19627: data = 8'hed;
      17'd19628: data = 8'hed;
      17'd19629: data = 8'hec;
      17'd19630: data = 8'heb;
      17'd19631: data = 8'heb;
      17'd19632: data = 8'heb;
      17'd19633: data = 8'heb;
      17'd19634: data = 8'he9;
      17'd19635: data = 8'heb;
      17'd19636: data = 8'he9;
      17'd19637: data = 8'he5;
      17'd19638: data = 8'he9;
      17'd19639: data = 8'heb;
      17'd19640: data = 8'he7;
      17'd19641: data = 8'he7;
      17'd19642: data = 8'he9;
      17'd19643: data = 8'heb;
      17'd19644: data = 8'heb;
      17'd19645: data = 8'he9;
      17'd19646: data = 8'he7;
      17'd19647: data = 8'he9;
      17'd19648: data = 8'hed;
      17'd19649: data = 8'hf1;
      17'd19650: data = 8'heb;
      17'd19651: data = 8'he3;
      17'd19652: data = 8'hdc;
      17'd19653: data = 8'hd8;
      17'd19654: data = 8'hdc;
      17'd19655: data = 8'hec;
      17'd19656: data = 8'hfc;
      17'd19657: data = 8'h02;
      17'd19658: data = 8'h01;
      17'd19659: data = 8'hfe;
      17'd19660: data = 8'h00;
      17'd19661: data = 8'hfa;
      17'd19662: data = 8'hf9;
      17'd19663: data = 8'hf1;
      17'd19664: data = 8'he3;
      17'd19665: data = 8'hdc;
      17'd19666: data = 8'he2;
      17'd19667: data = 8'hec;
      17'd19668: data = 8'hfa;
      17'd19669: data = 8'h09;
      17'd19670: data = 8'h0e;
      17'd19671: data = 8'h13;
      17'd19672: data = 8'h19;
      17'd19673: data = 8'h11;
      17'd19674: data = 8'h01;
      17'd19675: data = 8'hfd;
      17'd19676: data = 8'hfc;
      17'd19677: data = 8'h00;
      17'd19678: data = 8'h02;
      17'd19679: data = 8'hfe;
      17'd19680: data = 8'hf9;
      17'd19681: data = 8'hfd;
      17'd19682: data = 8'h06;
      17'd19683: data = 8'h11;
      17'd19684: data = 8'h23;
      17'd19685: data = 8'h31;
      17'd19686: data = 8'h33;
      17'd19687: data = 8'h29;
      17'd19688: data = 8'h13;
      17'd19689: data = 8'hfd;
      17'd19690: data = 8'hf1;
      17'd19691: data = 8'hf1;
      17'd19692: data = 8'hfd;
      17'd19693: data = 8'h13;
      17'd19694: data = 8'h29;
      17'd19695: data = 8'h35;
      17'd19696: data = 8'h35;
      17'd19697: data = 8'h2f;
      17'd19698: data = 8'h1f;
      17'd19699: data = 8'h15;
      17'd19700: data = 8'h0e;
      17'd19701: data = 8'h06;
      17'd19702: data = 8'h01;
      17'd19703: data = 8'h02;
      17'd19704: data = 8'h0a;
      17'd19705: data = 8'h0c;
      17'd19706: data = 8'h0e;
      17'd19707: data = 8'h12;
      17'd19708: data = 8'h1f;
      17'd19709: data = 8'h26;
      17'd19710: data = 8'h24;
      17'd19711: data = 8'h23;
      17'd19712: data = 8'h1a;
      17'd19713: data = 8'h16;
      17'd19714: data = 8'h11;
      17'd19715: data = 8'h04;
      17'd19716: data = 8'hfc;
      17'd19717: data = 8'hf4;
      17'd19718: data = 8'hf4;
      17'd19719: data = 8'hfc;
      17'd19720: data = 8'h01;
      17'd19721: data = 8'h05;
      17'd19722: data = 8'h0e;
      17'd19723: data = 8'h15;
      17'd19724: data = 8'h15;
      17'd19725: data = 8'h16;
      17'd19726: data = 8'h0e;
      17'd19727: data = 8'h06;
      17'd19728: data = 8'h02;
      17'd19729: data = 8'hfa;
      17'd19730: data = 8'hf5;
      17'd19731: data = 8'hf2;
      17'd19732: data = 8'hf2;
      17'd19733: data = 8'hf6;
      17'd19734: data = 8'h01;
      17'd19735: data = 8'h0a;
      17'd19736: data = 8'h12;
      17'd19737: data = 8'h1a;
      17'd19738: data = 8'h1e;
      17'd19739: data = 8'h1c;
      17'd19740: data = 8'h13;
      17'd19741: data = 8'h06;
      17'd19742: data = 8'hfd;
      17'd19743: data = 8'hf9;
      17'd19744: data = 8'hf9;
      17'd19745: data = 8'hfc;
      17'd19746: data = 8'h04;
      17'd19747: data = 8'h0c;
      17'd19748: data = 8'h0c;
      17'd19749: data = 8'h13;
      17'd19750: data = 8'h1a;
      17'd19751: data = 8'h19;
      17'd19752: data = 8'h19;
      17'd19753: data = 8'h16;
      17'd19754: data = 8'h0e;
      17'd19755: data = 8'h09;
      17'd19756: data = 8'h05;
      17'd19757: data = 8'h00;
      17'd19758: data = 8'hfd;
      17'd19759: data = 8'hfe;
      17'd19760: data = 8'h00;
      17'd19761: data = 8'h02;
      17'd19762: data = 8'h05;
      17'd19763: data = 8'h09;
      17'd19764: data = 8'h0e;
      17'd19765: data = 8'h0c;
      17'd19766: data = 8'h09;
      17'd19767: data = 8'h00;
      17'd19768: data = 8'hf6;
      17'd19769: data = 8'hef;
      17'd19770: data = 8'he7;
      17'd19771: data = 8'he7;
      17'd19772: data = 8'he3;
      17'd19773: data = 8'he3;
      17'd19774: data = 8'he9;
      17'd19775: data = 8'hf1;
      17'd19776: data = 8'hf5;
      17'd19777: data = 8'hf6;
      17'd19778: data = 8'hf9;
      17'd19779: data = 8'hf9;
      17'd19780: data = 8'hf2;
      17'd19781: data = 8'hed;
      17'd19782: data = 8'he9;
      17'd19783: data = 8'he7;
      17'd19784: data = 8'he7;
      17'd19785: data = 8'he7;
      17'd19786: data = 8'hec;
      17'd19787: data = 8'hef;
      17'd19788: data = 8'hf6;
      17'd19789: data = 8'hfd;
      17'd19790: data = 8'h00;
      17'd19791: data = 8'h04;
      17'd19792: data = 8'h05;
      17'd19793: data = 8'h02;
      17'd19794: data = 8'hfe;
      17'd19795: data = 8'hfd;
      17'd19796: data = 8'hfd;
      17'd19797: data = 8'hfd;
      17'd19798: data = 8'hfd;
      17'd19799: data = 8'h02;
      17'd19800: data = 8'h05;
      17'd19801: data = 8'h0a;
      17'd19802: data = 8'h11;
      17'd19803: data = 8'h13;
      17'd19804: data = 8'h16;
      17'd19805: data = 8'h15;
      17'd19806: data = 8'h16;
      17'd19807: data = 8'h16;
      17'd19808: data = 8'h11;
      17'd19809: data = 8'h0d;
      17'd19810: data = 8'h0c;
      17'd19811: data = 8'h0a;
      17'd19812: data = 8'h0a;
      17'd19813: data = 8'h0a;
      17'd19814: data = 8'h0c;
      17'd19815: data = 8'h11;
      17'd19816: data = 8'h12;
      17'd19817: data = 8'h13;
      17'd19818: data = 8'h0e;
      17'd19819: data = 8'h0c;
      17'd19820: data = 8'h0c;
      17'd19821: data = 8'h0a;
      17'd19822: data = 8'h09;
      17'd19823: data = 8'h01;
      17'd19824: data = 8'hfd;
      17'd19825: data = 8'hfa;
      17'd19826: data = 8'hf9;
      17'd19827: data = 8'hfc;
      17'd19828: data = 8'hfe;
      17'd19829: data = 8'h01;
      17'd19830: data = 8'h02;
      17'd19831: data = 8'h01;
      17'd19832: data = 8'hfa;
      17'd19833: data = 8'hf4;
      17'd19834: data = 8'hef;
      17'd19835: data = 8'heb;
      17'd19836: data = 8'he4;
      17'd19837: data = 8'he4;
      17'd19838: data = 8'he7;
      17'd19839: data = 8'hec;
      17'd19840: data = 8'hf4;
      17'd19841: data = 8'hf9;
      17'd19842: data = 8'hf9;
      17'd19843: data = 8'hf4;
      17'd19844: data = 8'hef;
      17'd19845: data = 8'heb;
      17'd19846: data = 8'he0;
      17'd19847: data = 8'hdb;
      17'd19848: data = 8'he2;
      17'd19849: data = 8'he9;
      17'd19850: data = 8'hef;
      17'd19851: data = 8'hed;
      17'd19852: data = 8'hf2;
      17'd19853: data = 8'hf5;
      17'd19854: data = 8'hf1;
      17'd19855: data = 8'heb;
      17'd19856: data = 8'he7;
      17'd19857: data = 8'he9;
      17'd19858: data = 8'heb;
      17'd19859: data = 8'hec;
      17'd19860: data = 8'hec;
      17'd19861: data = 8'hed;
      17'd19862: data = 8'he9;
      17'd19863: data = 8'he7;
      17'd19864: data = 8'he7;
      17'd19865: data = 8'he7;
      17'd19866: data = 8'heb;
      17'd19867: data = 8'hec;
      17'd19868: data = 8'hf1;
      17'd19869: data = 8'hf2;
      17'd19870: data = 8'hed;
      17'd19871: data = 8'hec;
      17'd19872: data = 8'hed;
      17'd19873: data = 8'he4;
      17'd19874: data = 8'hde;
      17'd19875: data = 8'he2;
      17'd19876: data = 8'he4;
      17'd19877: data = 8'he5;
      17'd19878: data = 8'hec;
      17'd19879: data = 8'hf1;
      17'd19880: data = 8'hed;
      17'd19881: data = 8'he9;
      17'd19882: data = 8'he4;
      17'd19883: data = 8'he3;
      17'd19884: data = 8'he5;
      17'd19885: data = 8'he7;
      17'd19886: data = 8'he7;
      17'd19887: data = 8'he4;
      17'd19888: data = 8'he7;
      17'd19889: data = 8'he5;
      17'd19890: data = 8'he5;
      17'd19891: data = 8'he7;
      17'd19892: data = 8'he4;
      17'd19893: data = 8'hf4;
      17'd19894: data = 8'hfc;
      17'd19895: data = 8'hf6;
      17'd19896: data = 8'hf6;
      17'd19897: data = 8'heb;
      17'd19898: data = 8'he9;
      17'd19899: data = 8'hfc;
      17'd19900: data = 8'h01;
      17'd19901: data = 8'hfd;
      17'd19902: data = 8'hfe;
      17'd19903: data = 8'h04;
      17'd19904: data = 8'h01;
      17'd19905: data = 8'hf9;
      17'd19906: data = 8'h05;
      17'd19907: data = 8'h19;
      17'd19908: data = 8'h15;
      17'd19909: data = 8'h13;
      17'd19910: data = 8'h1f;
      17'd19911: data = 8'h13;
      17'd19912: data = 8'h00;
      17'd19913: data = 8'h0c;
      17'd19914: data = 8'h11;
      17'd19915: data = 8'h11;
      17'd19916: data = 8'h13;
      17'd19917: data = 8'h19;
      17'd19918: data = 8'h1b;
      17'd19919: data = 8'h1f;
      17'd19920: data = 8'h26;
      17'd19921: data = 8'h1c;
      17'd19922: data = 8'h13;
      17'd19923: data = 8'h1c;
      17'd19924: data = 8'h1b;
      17'd19925: data = 8'h15;
      17'd19926: data = 8'h19;
      17'd19927: data = 8'h19;
      17'd19928: data = 8'h19;
      17'd19929: data = 8'h1c;
      17'd19930: data = 8'h1c;
      17'd19931: data = 8'h16;
      17'd19932: data = 8'h19;
      17'd19933: data = 8'h16;
      17'd19934: data = 8'h16;
      17'd19935: data = 8'h15;
      17'd19936: data = 8'h0e;
      17'd19937: data = 8'h0c;
      17'd19938: data = 8'h0c;
      17'd19939: data = 8'h0e;
      17'd19940: data = 8'h11;
      17'd19941: data = 8'h0a;
      17'd19942: data = 8'h0c;
      17'd19943: data = 8'h15;
      17'd19944: data = 8'h11;
      17'd19945: data = 8'h0c;
      17'd19946: data = 8'h09;
      17'd19947: data = 8'h01;
      17'd19948: data = 8'hf9;
      17'd19949: data = 8'hf5;
      17'd19950: data = 8'hf1;
      17'd19951: data = 8'he4;
      17'd19952: data = 8'he2;
      17'd19953: data = 8'hec;
      17'd19954: data = 8'hfd;
      17'd19955: data = 8'h0c;
      17'd19956: data = 8'h1a;
      17'd19957: data = 8'h1e;
      17'd19958: data = 8'h1c;
      17'd19959: data = 8'h13;
      17'd19960: data = 8'h01;
      17'd19961: data = 8'hec;
      17'd19962: data = 8'he2;
      17'd19963: data = 8'he3;
      17'd19964: data = 8'heb;
      17'd19965: data = 8'hf6;
      17'd19966: data = 8'h02;
      17'd19967: data = 8'h12;
      17'd19968: data = 8'h23;
      17'd19969: data = 8'h26;
      17'd19970: data = 8'h1f;
      17'd19971: data = 8'h1b;
      17'd19972: data = 8'h19;
      17'd19973: data = 8'h0e;
      17'd19974: data = 8'h05;
      17'd19975: data = 8'hfe;
      17'd19976: data = 8'hfd;
      17'd19977: data = 8'hfe;
      17'd19978: data = 8'h05;
      17'd19979: data = 8'h0e;
      17'd19980: data = 8'h13;
      17'd19981: data = 8'h1b;
      17'd19982: data = 8'h23;
      17'd19983: data = 8'h26;
      17'd19984: data = 8'h1f;
      17'd19985: data = 8'h13;
      17'd19986: data = 8'h0d;
      17'd19987: data = 8'h0c;
      17'd19988: data = 8'h04;
      17'd19989: data = 8'hfe;
      17'd19990: data = 8'hf6;
      17'd19991: data = 8'hf6;
      17'd19992: data = 8'hfc;
      17'd19993: data = 8'hfd;
      17'd19994: data = 8'h00;
      17'd19995: data = 8'h02;
      17'd19996: data = 8'h04;
      17'd19997: data = 8'h04;
      17'd19998: data = 8'h00;
      17'd19999: data = 8'hfa;
      17'd20000: data = 8'hf1;
      17'd20001: data = 8'he4;
      17'd20002: data = 8'hde;
      17'd20003: data = 8'hdb;
      17'd20004: data = 8'hdc;
      17'd20005: data = 8'he0;
      17'd20006: data = 8'he3;
      17'd20007: data = 8'he9;
      17'd20008: data = 8'hed;
      17'd20009: data = 8'hf5;
      17'd20010: data = 8'hf4;
      17'd20011: data = 8'hf5;
      17'd20012: data = 8'hf6;
      17'd20013: data = 8'hf4;
      17'd20014: data = 8'hf1;
      17'd20015: data = 8'hed;
      17'd20016: data = 8'heb;
      17'd20017: data = 8'he9;
      17'd20018: data = 8'heb;
      17'd20019: data = 8'hf2;
      17'd20020: data = 8'hfc;
      17'd20021: data = 8'h02;
      17'd20022: data = 8'h0c;
      17'd20023: data = 8'h12;
      17'd20024: data = 8'h15;
      17'd20025: data = 8'h16;
      17'd20026: data = 8'h16;
      17'd20027: data = 8'h13;
      17'd20028: data = 8'h11;
      17'd20029: data = 8'h0e;
      17'd20030: data = 8'h0d;
      17'd20031: data = 8'h11;
      17'd20032: data = 8'h15;
      17'd20033: data = 8'h1b;
      17'd20034: data = 8'h22;
      17'd20035: data = 8'h26;
      17'd20036: data = 8'h2b;
      17'd20037: data = 8'h2f;
      17'd20038: data = 8'h31;
      17'd20039: data = 8'h2b;
      17'd20040: data = 8'h24;
      17'd20041: data = 8'h1e;
      17'd20042: data = 8'h1a;
      17'd20043: data = 8'h1a;
      17'd20044: data = 8'h15;
      17'd20045: data = 8'h13;
      17'd20046: data = 8'h13;
      17'd20047: data = 8'h13;
      17'd20048: data = 8'h1a;
      17'd20049: data = 8'h19;
      17'd20050: data = 8'h16;
      17'd20051: data = 8'h13;
      17'd20052: data = 8'h12;
      17'd20053: data = 8'h0e;
      17'd20054: data = 8'h05;
      17'd20055: data = 8'h02;
      17'd20056: data = 8'hfa;
      17'd20057: data = 8'hf5;
      17'd20058: data = 8'hf1;
      17'd20059: data = 8'hed;
      17'd20060: data = 8'hef;
      17'd20061: data = 8'hef;
      17'd20062: data = 8'hef;
      17'd20063: data = 8'hf2;
      17'd20064: data = 8'hf4;
      17'd20065: data = 8'hf4;
      17'd20066: data = 8'hf1;
      17'd20067: data = 8'hec;
      17'd20068: data = 8'he7;
      17'd20069: data = 8'hdb;
      17'd20070: data = 8'hd3;
      17'd20071: data = 8'hd2;
      17'd20072: data = 8'hd2;
      17'd20073: data = 8'hda;
      17'd20074: data = 8'hde;
      17'd20075: data = 8'he3;
      17'd20076: data = 8'he9;
      17'd20077: data = 8'hec;
      17'd20078: data = 8'hef;
      17'd20079: data = 8'hf4;
      17'd20080: data = 8'hf4;
      17'd20081: data = 8'hed;
      17'd20082: data = 8'he9;
      17'd20083: data = 8'he4;
      17'd20084: data = 8'he2;
      17'd20085: data = 8'he3;
      17'd20086: data = 8'he5;
      17'd20087: data = 8'he9;
      17'd20088: data = 8'hef;
      17'd20089: data = 8'hf5;
      17'd20090: data = 8'hfc;
      17'd20091: data = 8'hfc;
      17'd20092: data = 8'hfd;
      17'd20093: data = 8'hfd;
      17'd20094: data = 8'hfc;
      17'd20095: data = 8'hf9;
      17'd20096: data = 8'hf2;
      17'd20097: data = 8'hed;
      17'd20098: data = 8'he5;
      17'd20099: data = 8'he2;
      17'd20100: data = 8'he2;
      17'd20101: data = 8'heb;
      17'd20102: data = 8'hf4;
      17'd20103: data = 8'hf9;
      17'd20104: data = 8'hfc;
      17'd20105: data = 8'hfa;
      17'd20106: data = 8'hf5;
      17'd20107: data = 8'hf4;
      17'd20108: data = 8'hef;
      17'd20109: data = 8'he9;
      17'd20110: data = 8'he4;
      17'd20111: data = 8'he3;
      17'd20112: data = 8'he0;
      17'd20113: data = 8'he2;
      17'd20114: data = 8'he4;
      17'd20115: data = 8'he4;
      17'd20116: data = 8'he4;
      17'd20117: data = 8'he3;
      17'd20118: data = 8'he4;
      17'd20119: data = 8'he7;
      17'd20120: data = 8'he5;
      17'd20121: data = 8'he4;
      17'd20122: data = 8'he4;
      17'd20123: data = 8'he2;
      17'd20124: data = 8'he0;
      17'd20125: data = 8'hdc;
      17'd20126: data = 8'hde;
      17'd20127: data = 8'he0;
      17'd20128: data = 8'he0;
      17'd20129: data = 8'he9;
      17'd20130: data = 8'hed;
      17'd20131: data = 8'hf4;
      17'd20132: data = 8'hfd;
      17'd20133: data = 8'h00;
      17'd20134: data = 8'h02;
      17'd20135: data = 8'h00;
      17'd20136: data = 8'h02;
      17'd20137: data = 8'h05;
      17'd20138: data = 8'h04;
      17'd20139: data = 8'h04;
      17'd20140: data = 8'h09;
      17'd20141: data = 8'h0c;
      17'd20142: data = 8'h0c;
      17'd20143: data = 8'h13;
      17'd20144: data = 8'h1a;
      17'd20145: data = 8'h22;
      17'd20146: data = 8'h27;
      17'd20147: data = 8'h2b;
      17'd20148: data = 8'h26;
      17'd20149: data = 8'h24;
      17'd20150: data = 8'h26;
      17'd20151: data = 8'h1c;
      17'd20152: data = 8'h15;
      17'd20153: data = 8'h13;
      17'd20154: data = 8'h16;
      17'd20155: data = 8'h16;
      17'd20156: data = 8'h1a;
      17'd20157: data = 8'h1e;
      17'd20158: data = 8'h23;
      17'd20159: data = 8'h27;
      17'd20160: data = 8'h29;
      17'd20161: data = 8'h24;
      17'd20162: data = 8'h23;
      17'd20163: data = 8'h26;
      17'd20164: data = 8'h1e;
      17'd20165: data = 8'h0e;
      17'd20166: data = 8'h04;
      17'd20167: data = 8'h02;
      17'd20168: data = 8'hfd;
      17'd20169: data = 8'hfe;
      17'd20170: data = 8'h05;
      17'd20171: data = 8'h13;
      17'd20172: data = 8'h23;
      17'd20173: data = 8'h24;
      17'd20174: data = 8'h1b;
      17'd20175: data = 8'h09;
      17'd20176: data = 8'hed;
      17'd20177: data = 8'hd1;
      17'd20178: data = 8'hc0;
      17'd20179: data = 8'hc2;
      17'd20180: data = 8'hce;
      17'd20181: data = 8'he7;
      17'd20182: data = 8'h0c;
      17'd20183: data = 8'h23;
      17'd20184: data = 8'h33;
      17'd20185: data = 8'h34;
      17'd20186: data = 8'h26;
      17'd20187: data = 8'h0c;
      17'd20188: data = 8'hed;
      17'd20189: data = 8'he4;
      17'd20190: data = 8'hde;
      17'd20191: data = 8'hdb;
      17'd20192: data = 8'he4;
      17'd20193: data = 8'hfa;
      17'd20194: data = 8'h12;
      17'd20195: data = 8'h24;
      17'd20196: data = 8'h2d;
      17'd20197: data = 8'h34;
      17'd20198: data = 8'h36;
      17'd20199: data = 8'h31;
      17'd20200: data = 8'h1f;
      17'd20201: data = 8'h0a;
      17'd20202: data = 8'h00;
      17'd20203: data = 8'hfc;
      17'd20204: data = 8'h00;
      17'd20205: data = 8'h04;
      17'd20206: data = 8'h0d;
      17'd20207: data = 8'h16;
      17'd20208: data = 8'h1b;
      17'd20209: data = 8'h23;
      17'd20210: data = 8'h1e;
      17'd20211: data = 8'h19;
      17'd20212: data = 8'h1a;
      17'd20213: data = 8'h19;
      17'd20214: data = 8'h16;
      17'd20215: data = 8'h0d;
      17'd20216: data = 8'h02;
      17'd20217: data = 8'hfc;
      17'd20218: data = 8'hf4;
      17'd20219: data = 8'hec;
      17'd20220: data = 8'he3;
      17'd20221: data = 8'he4;
      17'd20222: data = 8'hec;
      17'd20223: data = 8'hed;
      17'd20224: data = 8'he9;
      17'd20225: data = 8'hec;
      17'd20226: data = 8'hed;
      17'd20227: data = 8'hed;
      17'd20228: data = 8'he9;
      17'd20229: data = 8'he4;
      17'd20230: data = 8'he3;
      17'd20231: data = 8'hd6;
      17'd20232: data = 8'hcb;
      17'd20233: data = 8'hc4;
      17'd20234: data = 8'hc2;
      17'd20235: data = 8'hc9;
      17'd20236: data = 8'hd6;
      17'd20237: data = 8'he5;
      17'd20238: data = 8'hf5;
      17'd20239: data = 8'hfe;
      17'd20240: data = 8'h02;
      17'd20241: data = 8'h01;
      17'd20242: data = 8'hfc;
      17'd20243: data = 8'hf6;
      17'd20244: data = 8'hf1;
      17'd20245: data = 8'hf2;
      17'd20246: data = 8'hf4;
      17'd20247: data = 8'hf6;
      17'd20248: data = 8'h00;
      17'd20249: data = 8'h0a;
      17'd20250: data = 8'h16;
      17'd20251: data = 8'h22;
      17'd20252: data = 8'h33;
      17'd20253: data = 8'h3c;
      17'd20254: data = 8'h3d;
      17'd20255: data = 8'h3a;
      17'd20256: data = 8'h31;
      17'd20257: data = 8'h2b;
      17'd20258: data = 8'h26;
      17'd20259: data = 8'h27;
      17'd20260: data = 8'h29;
      17'd20261: data = 8'h2d;
      17'd20262: data = 8'h39;
      17'd20263: data = 8'h3a;
      17'd20264: data = 8'h39;
      17'd20265: data = 8'h36;
      17'd20266: data = 8'h35;
      17'd20267: data = 8'h3a;
      17'd20268: data = 8'h3c;
      17'd20269: data = 8'h36;
      17'd20270: data = 8'h31;
      17'd20271: data = 8'h2d;
      17'd20272: data = 8'h23;
      17'd20273: data = 8'h19;
      17'd20274: data = 8'h0e;
      17'd20275: data = 8'h09;
      17'd20276: data = 8'h0a;
      17'd20277: data = 8'h09;
      17'd20278: data = 8'h09;
      17'd20279: data = 8'h06;
      17'd20280: data = 8'h01;
      17'd20281: data = 8'hfe;
      17'd20282: data = 8'h00;
      17'd20283: data = 8'hfd;
      17'd20284: data = 8'hf9;
      17'd20285: data = 8'hf6;
      17'd20286: data = 8'hf2;
      17'd20287: data = 8'he9;
      17'd20288: data = 8'hda;
      17'd20289: data = 8'hce;
      17'd20290: data = 8'hc9;
      17'd20291: data = 8'hc6;
      17'd20292: data = 8'hca;
      17'd20293: data = 8'hd5;
      17'd20294: data = 8'hde;
      17'd20295: data = 8'he3;
      17'd20296: data = 8'he9;
      17'd20297: data = 8'heb;
      17'd20298: data = 8'he7;
      17'd20299: data = 8'hde;
      17'd20300: data = 8'hce;
      17'd20301: data = 8'hc4;
      17'd20302: data = 8'hbd;
      17'd20303: data = 8'hc0;
      17'd20304: data = 8'hca;
      17'd20305: data = 8'hd6;
      17'd20306: data = 8'he5;
      17'd20307: data = 8'hf5;
      17'd20308: data = 8'h01;
      17'd20309: data = 8'h09;
      17'd20310: data = 8'h04;
      17'd20311: data = 8'hfc;
      17'd20312: data = 8'hf6;
      17'd20313: data = 8'hed;
      17'd20314: data = 8'he5;
      17'd20315: data = 8'he5;
      17'd20316: data = 8'hec;
      17'd20317: data = 8'hf2;
      17'd20318: data = 8'hf4;
      17'd20319: data = 8'hfa;
      17'd20320: data = 8'h01;
      17'd20321: data = 8'h05;
      17'd20322: data = 8'h06;
      17'd20323: data = 8'h06;
      17'd20324: data = 8'h02;
      17'd20325: data = 8'hfc;
      17'd20326: data = 8'hf6;
      17'd20327: data = 8'hf4;
      17'd20328: data = 8'heb;
      17'd20329: data = 8'he5;
      17'd20330: data = 8'he3;
      17'd20331: data = 8'he2;
      17'd20332: data = 8'he3;
      17'd20333: data = 8'he4;
      17'd20334: data = 8'he5;
      17'd20335: data = 8'he9;
      17'd20336: data = 8'hef;
      17'd20337: data = 8'hf1;
      17'd20338: data = 8'hf1;
      17'd20339: data = 8'hf1;
      17'd20340: data = 8'heb;
      17'd20341: data = 8'he4;
      17'd20342: data = 8'hd8;
      17'd20343: data = 8'hca;
      17'd20344: data = 8'hc5;
      17'd20345: data = 8'hc2;
      17'd20346: data = 8'hc4;
      17'd20347: data = 8'hc6;
      17'd20348: data = 8'hd5;
      17'd20349: data = 8'hde;
      17'd20350: data = 8'he2;
      17'd20351: data = 8'hec;
      17'd20352: data = 8'hf2;
      17'd20353: data = 8'hec;
      17'd20354: data = 8'he4;
      17'd20355: data = 8'hde;
      17'd20356: data = 8'hd6;
      17'd20357: data = 8'hd8;
      17'd20358: data = 8'hdc;
      17'd20359: data = 8'he7;
      17'd20360: data = 8'hf1;
      17'd20361: data = 8'hfe;
      17'd20362: data = 8'h0d;
      17'd20363: data = 8'h1c;
      17'd20364: data = 8'h23;
      17'd20365: data = 8'h23;
      17'd20366: data = 8'h22;
      17'd20367: data = 8'h1b;
      17'd20368: data = 8'h1a;
      17'd20369: data = 8'h13;
      17'd20370: data = 8'h15;
      17'd20371: data = 8'h16;
      17'd20372: data = 8'h1e;
      17'd20373: data = 8'h1f;
      17'd20374: data = 8'h23;
      17'd20375: data = 8'h2c;
      17'd20376: data = 8'h33;
      17'd20377: data = 8'h2f;
      17'd20378: data = 8'h29;
      17'd20379: data = 8'h31;
      17'd20380: data = 8'h29;
      17'd20381: data = 8'h29;
      17'd20382: data = 8'h2d;
      17'd20383: data = 8'h26;
      17'd20384: data = 8'h1f;
      17'd20385: data = 8'h19;
      17'd20386: data = 8'h13;
      17'd20387: data = 8'h0e;
      17'd20388: data = 8'h01;
      17'd20389: data = 8'h06;
      17'd20390: data = 8'h0c;
      17'd20391: data = 8'h11;
      17'd20392: data = 8'h1f;
      17'd20393: data = 8'h24;
      17'd20394: data = 8'h31;
      17'd20395: data = 8'h26;
      17'd20396: data = 8'h06;
      17'd20397: data = 8'hf6;
      17'd20398: data = 8'hd3;
      17'd20399: data = 8'hb3;
      17'd20400: data = 8'ha6;
      17'd20401: data = 8'ha8;
      17'd20402: data = 8'hc0;
      17'd20403: data = 8'hda;
      17'd20404: data = 8'h12;
      17'd20405: data = 8'h35;
      17'd20406: data = 8'h3e;
      17'd20407: data = 8'h47;
      17'd20408: data = 8'h33;
      17'd20409: data = 8'h12;
      17'd20410: data = 8'hf1;
      17'd20411: data = 8'hd8;
      17'd20412: data = 8'hcd;
      17'd20413: data = 8'hc5;
      17'd20414: data = 8'hcd;
      17'd20415: data = 8'he3;
      17'd20416: data = 8'h00;
      17'd20417: data = 8'h22;
      17'd20418: data = 8'h3c;
      17'd20419: data = 8'h4d;
      17'd20420: data = 8'h56;
      17'd20421: data = 8'h4d;
      17'd20422: data = 8'h3d;
      17'd20423: data = 8'h26;
      17'd20424: data = 8'h0d;
      17'd20425: data = 8'h00;
      17'd20426: data = 8'hfc;
      17'd20427: data = 8'h00;
      17'd20428: data = 8'h09;
      17'd20429: data = 8'h11;
      17'd20430: data = 8'h1b;
      17'd20431: data = 8'h1c;
      17'd20432: data = 8'h1b;
      17'd20433: data = 8'h24;
      17'd20434: data = 8'h2b;
      17'd20435: data = 8'h2d;
      17'd20436: data = 8'h2f;
      17'd20437: data = 8'h2b;
      17'd20438: data = 8'h1a;
      17'd20439: data = 8'h04;
      17'd20440: data = 8'hfa;
      17'd20441: data = 8'heb;
      17'd20442: data = 8'hd6;
      17'd20443: data = 8'hd3;
      17'd20444: data = 8'hd1;
      17'd20445: data = 8'hcb;
      17'd20446: data = 8'hc9;
      17'd20447: data = 8'hd1;
      17'd20448: data = 8'hdc;
      17'd20449: data = 8'heb;
      17'd20450: data = 8'hf6;
      17'd20451: data = 8'hfc;
      17'd20452: data = 8'hf9;
      17'd20453: data = 8'he5;
      17'd20454: data = 8'hc6;
      17'd20455: data = 8'hb0;
      17'd20456: data = 8'ha3;
      17'd20457: data = 8'h9b;
      17'd20458: data = 8'ha6;
      17'd20459: data = 8'hbd;
      17'd20460: data = 8'hd2;
      17'd20461: data = 8'he2;
      17'd20462: data = 8'hf5;
      17'd20463: data = 8'h06;
      17'd20464: data = 8'h0e;
      17'd20465: data = 8'h12;
      17'd20466: data = 8'h13;
      17'd20467: data = 8'h0d;
      17'd20468: data = 8'h00;
      17'd20469: data = 8'hf6;
      17'd20470: data = 8'hf2;
      17'd20471: data = 8'hf1;
      17'd20472: data = 8'hfc;
      17'd20473: data = 8'h0e;
      17'd20474: data = 8'h26;
      17'd20475: data = 8'h3c;
      17'd20476: data = 8'h47;
      17'd20477: data = 8'h4d;
      17'd20478: data = 8'h4e;
      17'd20479: data = 8'h52;
      17'd20480: data = 8'h52;
      17'd20481: data = 8'h52;
      17'd20482: data = 8'h53;
      17'd20483: data = 8'h4e;
      17'd20484: data = 8'h45;
      17'd20485: data = 8'h3e;
      17'd20486: data = 8'h35;
      17'd20487: data = 8'h2d;
      17'd20488: data = 8'h31;
      17'd20489: data = 8'h3a;
      17'd20490: data = 8'h43;
      17'd20491: data = 8'h42;
      17'd20492: data = 8'h43;
      17'd20493: data = 8'h42;
      17'd20494: data = 8'h39;
      17'd20495: data = 8'h36;
      17'd20496: data = 8'h2f;
      17'd20497: data = 8'h22;
      17'd20498: data = 8'h19;
      17'd20499: data = 8'h05;
      17'd20500: data = 8'hf2;
      17'd20501: data = 8'he5;
      17'd20502: data = 8'hde;
      17'd20503: data = 8'hdc;
      17'd20504: data = 8'he2;
      17'd20505: data = 8'hec;
      17'd20506: data = 8'hf6;
      17'd20507: data = 8'h01;
      17'd20508: data = 8'h04;
      17'd20509: data = 8'hf4;
      17'd20510: data = 8'hda;
      17'd20511: data = 8'hcb;
      17'd20512: data = 8'hc2;
      17'd20513: data = 8'hb3;
      17'd20514: data = 8'hbb;
      17'd20515: data = 8'hbd;
      17'd20516: data = 8'hc2;
      17'd20517: data = 8'hce;
      17'd20518: data = 8'hda;
      17'd20519: data = 8'he2;
      17'd20520: data = 8'hdc;
      17'd20521: data = 8'he2;
      17'd20522: data = 8'he2;
      17'd20523: data = 8'hda;
      17'd20524: data = 8'hdb;
      17'd20525: data = 8'hd6;
      17'd20526: data = 8'hda;
      17'd20527: data = 8'he2;
      17'd20528: data = 8'he5;
      17'd20529: data = 8'heb;
      17'd20530: data = 8'hfc;
      17'd20531: data = 8'h09;
      17'd20532: data = 8'h00;
      17'd20533: data = 8'hfe;
      17'd20534: data = 8'h02;
      17'd20535: data = 8'hfd;
      17'd20536: data = 8'h02;
      17'd20537: data = 8'h0d;
      17'd20538: data = 8'h19;
      17'd20539: data = 8'h13;
      17'd20540: data = 8'h11;
      17'd20541: data = 8'h09;
      17'd20542: data = 8'hfe;
      17'd20543: data = 8'h00;
      17'd20544: data = 8'hfa;
      17'd20545: data = 8'hf5;
      17'd20546: data = 8'hf2;
      17'd20547: data = 8'hf4;
      17'd20548: data = 8'hf6;
      17'd20549: data = 8'hf4;
      17'd20550: data = 8'hfe;
      17'd20551: data = 8'hf9;
      17'd20552: data = 8'hf1;
      17'd20553: data = 8'hf1;
      17'd20554: data = 8'he5;
      17'd20555: data = 8'hdb;
      17'd20556: data = 8'hcb;
      17'd20557: data = 8'hc5;
      17'd20558: data = 8'hc2;
      17'd20559: data = 8'hc4;
      17'd20560: data = 8'hce;
      17'd20561: data = 8'hce;
      17'd20562: data = 8'hd8;
      17'd20563: data = 8'hda;
      17'd20564: data = 8'hcb;
      17'd20565: data = 8'hc5;
      17'd20566: data = 8'hc6;
      17'd20567: data = 8'hc4;
      17'd20568: data = 8'hbc;
      17'd20569: data = 8'hc5;
      17'd20570: data = 8'hca;
      17'd20571: data = 8'hc6;
      17'd20572: data = 8'hd3;
      17'd20573: data = 8'hda;
      17'd20574: data = 8'hd8;
      17'd20575: data = 8'hdb;
      17'd20576: data = 8'hde;
      17'd20577: data = 8'hde;
      17'd20578: data = 8'he4;
      17'd20579: data = 8'hed;
      17'd20580: data = 8'hf2;
      17'd20581: data = 8'hfe;
      17'd20582: data = 8'h0a;
      17'd20583: data = 8'h13;
      17'd20584: data = 8'h22;
      17'd20585: data = 8'h27;
      17'd20586: data = 8'h26;
      17'd20587: data = 8'h1e;
      17'd20588: data = 8'h1c;
      17'd20589: data = 8'h1b;
      17'd20590: data = 8'h1c;
      17'd20591: data = 8'h27;
      17'd20592: data = 8'h31;
      17'd20593: data = 8'h33;
      17'd20594: data = 8'h3a;
      17'd20595: data = 8'h3d;
      17'd20596: data = 8'h3a;
      17'd20597: data = 8'h3a;
      17'd20598: data = 8'h33;
      17'd20599: data = 8'h33;
      17'd20600: data = 8'h2f;
      17'd20601: data = 8'h2b;
      17'd20602: data = 8'h26;
      17'd20603: data = 8'h22;
      17'd20604: data = 8'h1c;
      17'd20605: data = 8'h12;
      17'd20606: data = 8'h11;
      17'd20607: data = 8'h1e;
      17'd20608: data = 8'h19;
      17'd20609: data = 8'h16;
      17'd20610: data = 8'h16;
      17'd20611: data = 8'h0d;
      17'd20612: data = 8'h0c;
      17'd20613: data = 8'h0e;
      17'd20614: data = 8'h0c;
      17'd20615: data = 8'hfc;
      17'd20616: data = 8'hf6;
      17'd20617: data = 8'hd8;
      17'd20618: data = 8'hb4;
      17'd20619: data = 8'haa;
      17'd20620: data = 8'hab;
      17'd20621: data = 8'hb4;
      17'd20622: data = 8'hc9;
      17'd20623: data = 8'hf9;
      17'd20624: data = 8'h16;
      17'd20625: data = 8'h22;
      17'd20626: data = 8'h31;
      17'd20627: data = 8'h2b;
      17'd20628: data = 8'h12;
      17'd20629: data = 8'h00;
      17'd20630: data = 8'hf5;
      17'd20631: data = 8'he4;
      17'd20632: data = 8'hdb;
      17'd20633: data = 8'hdb;
      17'd20634: data = 8'hd6;
      17'd20635: data = 8'he7;
      17'd20636: data = 8'h05;
      17'd20637: data = 8'h24;
      17'd20638: data = 8'h3c;
      17'd20639: data = 8'h56;
      17'd20640: data = 8'h60;
      17'd20641: data = 8'h4d;
      17'd20642: data = 8'h3d;
      17'd20643: data = 8'h31;
      17'd20644: data = 8'h1f;
      17'd20645: data = 8'h15;
      17'd20646: data = 8'h1b;
      17'd20647: data = 8'h1b;
      17'd20648: data = 8'h11;
      17'd20649: data = 8'h12;
      17'd20650: data = 8'h0a;
      17'd20651: data = 8'h05;
      17'd20652: data = 8'h12;
      17'd20653: data = 8'h1e;
      17'd20654: data = 8'h24;
      17'd20655: data = 8'h2d;
      17'd20656: data = 8'h2b;
      17'd20657: data = 8'h1a;
      17'd20658: data = 8'h0d;
      17'd20659: data = 8'h02;
      17'd20660: data = 8'hf2;
      17'd20661: data = 8'he5;
      17'd20662: data = 8'hde;
      17'd20663: data = 8'hc5;
      17'd20664: data = 8'hb0;
      17'd20665: data = 8'ha4;
      17'd20666: data = 8'ha1;
      17'd20667: data = 8'ha6;
      17'd20668: data = 8'hbd;
      17'd20669: data = 8'hd8;
      17'd20670: data = 8'he3;
      17'd20671: data = 8'heb;
      17'd20672: data = 8'hec;
      17'd20673: data = 8'hdc;
      17'd20674: data = 8'hcb;
      17'd20675: data = 8'hc2;
      17'd20676: data = 8'hb3;
      17'd20677: data = 8'hb1;
      17'd20678: data = 8'hb3;
      17'd20679: data = 8'hb4;
      17'd20680: data = 8'hbb;
      17'd20681: data = 8'hc9;
      17'd20682: data = 8'hdc;
      17'd20683: data = 8'hef;
      17'd20684: data = 8'h11;
      17'd20685: data = 8'h26;
      17'd20686: data = 8'h31;
      17'd20687: data = 8'h2f;
      17'd20688: data = 8'h29;
      17'd20689: data = 8'h23;
      17'd20690: data = 8'h1a;
      17'd20691: data = 8'h1f;
      17'd20692: data = 8'h2b;
      17'd20693: data = 8'h2f;
      17'd20694: data = 8'h34;
      17'd20695: data = 8'h3c;
      17'd20696: data = 8'h3d;
      17'd20697: data = 8'h40;
      17'd20698: data = 8'h4e;
      17'd20699: data = 8'h57;
      17'd20700: data = 8'h64;
      17'd20701: data = 8'h6d;
      17'd20702: data = 8'h6a;
      17'd20703: data = 8'h65;
      17'd20704: data = 8'h63;
      17'd20705: data = 8'h56;
      17'd20706: data = 8'h4a;
      17'd20707: data = 8'h47;
      17'd20708: data = 8'h3e;
      17'd20709: data = 8'h31;
      17'd20710: data = 8'h24;
      17'd20711: data = 8'h1b;
      17'd20712: data = 8'h0d;
      17'd20713: data = 8'h0d;
      17'd20714: data = 8'h16;
      17'd20715: data = 8'h19;
      17'd20716: data = 8'h22;
      17'd20717: data = 8'h23;
      17'd20718: data = 8'h13;
      17'd20719: data = 8'h01;
      17'd20720: data = 8'hf4;
      17'd20721: data = 8'he4;
      17'd20722: data = 8'hd6;
      17'd20723: data = 8'hce;
      17'd20724: data = 8'hc6;
      17'd20725: data = 8'hc1;
      17'd20726: data = 8'hbd;
      17'd20727: data = 8'hc0;
      17'd20728: data = 8'hc1;
      17'd20729: data = 8'hd1;
      17'd20730: data = 8'hdc;
      17'd20731: data = 8'he0;
      17'd20732: data = 8'he5;
      17'd20733: data = 8'he4;
      17'd20734: data = 8'hd6;
      17'd20735: data = 8'hcd;
      17'd20736: data = 8'hca;
      17'd20737: data = 8'hca;
      17'd20738: data = 8'hce;
      17'd20739: data = 8'hd8;
      17'd20740: data = 8'hde;
      17'd20741: data = 8'he5;
      17'd20742: data = 8'he9;
      17'd20743: data = 8'hef;
      17'd20744: data = 8'hfa;
      17'd20745: data = 8'h01;
      17'd20746: data = 8'h12;
      17'd20747: data = 8'h15;
      17'd20748: data = 8'h1a;
      17'd20749: data = 8'h15;
      17'd20750: data = 8'h13;
      17'd20751: data = 8'h13;
      17'd20752: data = 8'h13;
      17'd20753: data = 8'h15;
      17'd20754: data = 8'h0e;
      17'd20755: data = 8'h11;
      17'd20756: data = 8'h0c;
      17'd20757: data = 8'h0c;
      17'd20758: data = 8'h0c;
      17'd20759: data = 8'h0d;
      17'd20760: data = 8'h0a;
      17'd20761: data = 8'h0a;
      17'd20762: data = 8'h12;
      17'd20763: data = 8'h0d;
      17'd20764: data = 8'h02;
      17'd20765: data = 8'hfc;
      17'd20766: data = 8'hed;
      17'd20767: data = 8'hdc;
      17'd20768: data = 8'hd3;
      17'd20769: data = 8'hcd;
      17'd20770: data = 8'hd3;
      17'd20771: data = 8'hce;
      17'd20772: data = 8'hbb;
      17'd20773: data = 8'hd5;
      17'd20774: data = 8'h04;
      17'd20775: data = 8'hd8;
      17'd20776: data = 8'ha1;
      17'd20777: data = 8'hcb;
      17'd20778: data = 8'he0;
      17'd20779: data = 8'hc1;
      17'd20780: data = 8'hbc;
      17'd20781: data = 8'hb3;
      17'd20782: data = 8'hb3;
      17'd20783: data = 8'hb3;
      17'd20784: data = 8'hab;
      17'd20785: data = 8'hb1;
      17'd20786: data = 8'hbd;
      17'd20787: data = 8'hc4;
      17'd20788: data = 8'hc1;
      17'd20789: data = 8'hcb;
      17'd20790: data = 8'hd6;
      17'd20791: data = 8'hde;
      17'd20792: data = 8'he7;
      17'd20793: data = 8'hec;
      17'd20794: data = 8'heb;
      17'd20795: data = 8'hf1;
      17'd20796: data = 8'hfa;
      17'd20797: data = 8'hf9;
      17'd20798: data = 8'h02;
      17'd20799: data = 8'h09;
      17'd20800: data = 8'h16;
      17'd20801: data = 8'h23;
      17'd20802: data = 8'h22;
      17'd20803: data = 8'h2d;
      17'd20804: data = 8'h31;
      17'd20805: data = 8'h34;
      17'd20806: data = 8'h3a;
      17'd20807: data = 8'h2c;
      17'd20808: data = 8'h2f;
      17'd20809: data = 8'h31;
      17'd20810: data = 8'h27;
      17'd20811: data = 8'h34;
      17'd20812: data = 8'h35;
      17'd20813: data = 8'h33;
      17'd20814: data = 8'h2d;
      17'd20815: data = 8'h35;
      17'd20816: data = 8'h39;
      17'd20817: data = 8'h27;
      17'd20818: data = 8'h2b;
      17'd20819: data = 8'h29;
      17'd20820: data = 8'h1a;
      17'd20821: data = 8'h13;
      17'd20822: data = 8'h05;
      17'd20823: data = 8'hfe;
      17'd20824: data = 8'h02;
      17'd20825: data = 8'h04;
      17'd20826: data = 8'hfd;
      17'd20827: data = 8'h05;
      17'd20828: data = 8'h01;
      17'd20829: data = 8'h09;
      17'd20830: data = 8'h0c;
      17'd20831: data = 8'h0c;
      17'd20832: data = 8'h0e;
      17'd20833: data = 8'hf5;
      17'd20834: data = 8'he9;
      17'd20835: data = 8'hc9;
      17'd20836: data = 8'hab;
      17'd20837: data = 8'ha1;
      17'd20838: data = 8'h9d;
      17'd20839: data = 8'ha8;
      17'd20840: data = 8'hc2;
      17'd20841: data = 8'hed;
      17'd20842: data = 8'h0c;
      17'd20843: data = 8'h1c;
      17'd20844: data = 8'h31;
      17'd20845: data = 8'h3e;
      17'd20846: data = 8'h2f;
      17'd20847: data = 8'h1e;
      17'd20848: data = 8'h15;
      17'd20849: data = 8'hfa;
      17'd20850: data = 8'hec;
      17'd20851: data = 8'hec;
      17'd20852: data = 8'hec;
      17'd20853: data = 8'hf5;
      17'd20854: data = 8'h11;
      17'd20855: data = 8'h24;
      17'd20856: data = 8'h31;
      17'd20857: data = 8'h4a;
      17'd20858: data = 8'h56;
      17'd20859: data = 8'h54;
      17'd20860: data = 8'h56;
      17'd20861: data = 8'h4a;
      17'd20862: data = 8'h3e;
      17'd20863: data = 8'h39;
      17'd20864: data = 8'h33;
      17'd20865: data = 8'h2d;
      17'd20866: data = 8'h23;
      17'd20867: data = 8'h1a;
      17'd20868: data = 8'h05;
      17'd20869: data = 8'hf6;
      17'd20870: data = 8'hf6;
      17'd20871: data = 8'hf6;
      17'd20872: data = 8'hf6;
      17'd20873: data = 8'h00;
      17'd20874: data = 8'h02;
      17'd20875: data = 8'h00;
      17'd20876: data = 8'hfe;
      17'd20877: data = 8'h04;
      17'd20878: data = 8'h01;
      17'd20879: data = 8'hed;
      17'd20880: data = 8'he2;
      17'd20881: data = 8'hce;
      17'd20882: data = 8'hac;
      17'd20883: data = 8'h9a;
      17'd20884: data = 8'h8c;
      17'd20885: data = 8'h83;
      17'd20886: data = 8'h89;
      17'd20887: data = 8'h94;
      17'd20888: data = 8'ha8;
      17'd20889: data = 8'hbc;
      17'd20890: data = 8'hcd;
      17'd20891: data = 8'hd3;
      17'd20892: data = 8'hd5;
      17'd20893: data = 8'hdc;
      17'd20894: data = 8'hd8;
      17'd20895: data = 8'hd8;
      17'd20896: data = 8'hd8;
      17'd20897: data = 8'hd2;
      17'd20898: data = 8'hcd;
      17'd20899: data = 8'hce;
      17'd20900: data = 8'hd3;
      17'd20901: data = 8'he2;
      17'd20902: data = 8'hfd;
      17'd20903: data = 8'h16;
      17'd20904: data = 8'h23;
      17'd20905: data = 8'h2f;
      17'd20906: data = 8'h3a;
      17'd20907: data = 8'h3d;
      17'd20908: data = 8'h43;
      17'd20909: data = 8'h52;
      17'd20910: data = 8'h5c;
      17'd20911: data = 8'h64;
      17'd20912: data = 8'h6d;
      17'd20913: data = 8'h6a;
      17'd20914: data = 8'h5b;
      17'd20915: data = 8'h4a;
      17'd20916: data = 8'h46;
      17'd20917: data = 8'h46;
      17'd20918: data = 8'h4e;
      17'd20919: data = 8'h4f;
      17'd20920: data = 8'h4d;
      17'd20921: data = 8'h4a;
      17'd20922: data = 8'h46;
      17'd20923: data = 8'h46;
      17'd20924: data = 8'h4d;
      17'd20925: data = 8'h56;
      17'd20926: data = 8'h56;
      17'd20927: data = 8'h46;
      17'd20928: data = 8'h34;
      17'd20929: data = 8'h1b;
      17'd20930: data = 8'hfe;
      17'd20931: data = 8'he9;
      17'd20932: data = 8'he2;
      17'd20933: data = 8'hdb;
      17'd20934: data = 8'hda;
      17'd20935: data = 8'hda;
      17'd20936: data = 8'hd6;
      17'd20937: data = 8'hd6;
      17'd20938: data = 8'hda;
      17'd20939: data = 8'hdc;
      17'd20940: data = 8'he3;
      17'd20941: data = 8'he5;
      17'd20942: data = 8'hde;
      17'd20943: data = 8'hd3;
      17'd20944: data = 8'hcd;
      17'd20945: data = 8'hc1;
      17'd20946: data = 8'hc0;
      17'd20947: data = 8'hc5;
      17'd20948: data = 8'hca;
      17'd20949: data = 8'hd3;
      17'd20950: data = 8'hda;
      17'd20951: data = 8'hdb;
      17'd20952: data = 8'hd8;
      17'd20953: data = 8'he0;
      17'd20954: data = 8'he5;
      17'd20955: data = 8'hed;
      17'd20956: data = 8'hfc;
      17'd20957: data = 8'h0d;
      17'd20958: data = 8'h13;
      17'd20959: data = 8'h12;
      17'd20960: data = 8'h1b;
      17'd20961: data = 8'h1f;
      17'd20962: data = 8'h24;
      17'd20963: data = 8'h26;
      17'd20964: data = 8'h2b;
      17'd20965: data = 8'h27;
      17'd20966: data = 8'h26;
      17'd20967: data = 8'h24;
      17'd20968: data = 8'h1c;
      17'd20969: data = 8'h1f;
      17'd20970: data = 8'h24;
      17'd20971: data = 8'h27;
      17'd20972: data = 8'h2b;
      17'd20973: data = 8'h2d;
      17'd20974: data = 8'h26;
      17'd20975: data = 8'h1c;
      17'd20976: data = 8'h13;
      17'd20977: data = 8'h06;
      17'd20978: data = 8'hfd;
      17'd20979: data = 8'hf6;
      17'd20980: data = 8'hf1;
      17'd20981: data = 8'he5;
      17'd20982: data = 8'hde;
      17'd20983: data = 8'hd6;
      17'd20984: data = 8'hcd;
      17'd20985: data = 8'hca;
      17'd20986: data = 8'hc9;
      17'd20987: data = 8'hc2;
      17'd20988: data = 8'hc2;
      17'd20989: data = 8'hc2;
      17'd20990: data = 8'hbd;
      17'd20991: data = 8'hbb;
      17'd20992: data = 8'hb5;
      17'd20993: data = 8'hb8;
      17'd20994: data = 8'hbb;
      17'd20995: data = 8'hbd;
      17'd20996: data = 8'hc0;
      17'd20997: data = 8'hc0;
      17'd20998: data = 8'hbc;
      17'd20999: data = 8'hb8;
      17'd21000: data = 8'hb3;
      17'd21001: data = 8'hb4;
      17'd21002: data = 8'hb9;
      17'd21003: data = 8'hc1;
      17'd21004: data = 8'hc6;
      17'd21005: data = 8'hd1;
      17'd21006: data = 8'hdc;
      17'd21007: data = 8'he9;
      17'd21008: data = 8'hf5;
      17'd21009: data = 8'hfe;
      17'd21010: data = 8'h02;
      17'd21011: data = 8'h0a;
      17'd21012: data = 8'h0a;
      17'd21013: data = 8'h06;
      17'd21014: data = 8'h0a;
      17'd21015: data = 8'h0a;
      17'd21016: data = 8'h11;
      17'd21017: data = 8'h1e;
      17'd21018: data = 8'h23;
      17'd21019: data = 8'h29;
      17'd21020: data = 8'h33;
      17'd21021: data = 8'h35;
      17'd21022: data = 8'h3a;
      17'd21023: data = 8'h3e;
      17'd21024: data = 8'h3d;
      17'd21025: data = 8'h43;
      17'd21026: data = 8'h40;
      17'd21027: data = 8'h31;
      17'd21028: data = 8'h31;
      17'd21029: data = 8'h24;
      17'd21030: data = 8'h1f;
      17'd21031: data = 8'h1b;
      17'd21032: data = 8'h16;
      17'd21033: data = 8'h15;
      17'd21034: data = 8'h0c;
      17'd21035: data = 8'h0d;
      17'd21036: data = 8'h02;
      17'd21037: data = 8'h02;
      17'd21038: data = 8'h06;
      17'd21039: data = 8'hfc;
      17'd21040: data = 8'hf4;
      17'd21041: data = 8'h04;
      17'd21042: data = 8'hf5;
      17'd21043: data = 8'hf1;
      17'd21044: data = 8'hf6;
      17'd21045: data = 8'hec;
      17'd21046: data = 8'he4;
      17'd21047: data = 8'he3;
      17'd21048: data = 8'he5;
      17'd21049: data = 8'heb;
      17'd21050: data = 8'hf9;
      17'd21051: data = 8'hf4;
      17'd21052: data = 8'hf4;
      17'd21053: data = 8'heb;
      17'd21054: data = 8'hd3;
      17'd21055: data = 8'hc1;
      17'd21056: data = 8'hb5;
      17'd21057: data = 8'hb9;
      17'd21058: data = 8'hb9;
      17'd21059: data = 8'hd2;
      17'd21060: data = 8'hfa;
      17'd21061: data = 8'h0e;
      17'd21062: data = 8'h22;
      17'd21063: data = 8'h40;
      17'd21064: data = 8'h4a;
      17'd21065: data = 8'h4d;
      17'd21066: data = 8'h4f;
      17'd21067: data = 8'h4a;
      17'd21068: data = 8'h35;
      17'd21069: data = 8'h1c;
      17'd21070: data = 8'h15;
      17'd21071: data = 8'h04;
      17'd21072: data = 8'h06;
      17'd21073: data = 8'h1a;
      17'd21074: data = 8'h2c;
      17'd21075: data = 8'h3a;
      17'd21076: data = 8'h46;
      17'd21077: data = 8'h53;
      17'd21078: data = 8'h4e;
      17'd21079: data = 8'h43;
      17'd21080: data = 8'h45;
      17'd21081: data = 8'h42;
      17'd21082: data = 8'h3d;
      17'd21083: data = 8'h34;
      17'd21084: data = 8'h26;
      17'd21085: data = 8'h1b;
      17'd21086: data = 8'h04;
      17'd21087: data = 8'hf1;
      17'd21088: data = 8'heb;
      17'd21089: data = 8'hf1;
      17'd21090: data = 8'he3;
      17'd21091: data = 8'hce;
      17'd21092: data = 8'hce;
      17'd21093: data = 8'hca;
      17'd21094: data = 8'hc1;
      17'd21095: data = 8'hc5;
      17'd21096: data = 8'hd2;
      17'd21097: data = 8'hd5;
      17'd21098: data = 8'hdb;
      17'd21099: data = 8'he2;
      17'd21100: data = 8'hd3;
      17'd21101: data = 8'hc0;
      17'd21102: data = 8'hae;
      17'd21103: data = 8'h9a;
      17'd21104: data = 8'h90;
      17'd21105: data = 8'h8a;
      17'd21106: data = 8'h8d;
      17'd21107: data = 8'h94;
      17'd21108: data = 8'h9d;
      17'd21109: data = 8'ha6;
      17'd21110: data = 8'hb8;
      17'd21111: data = 8'hcb;
      17'd21112: data = 8'he4;
      17'd21113: data = 8'hf9;
      17'd21114: data = 8'h04;
      17'd21115: data = 8'h09;
      17'd21116: data = 8'h00;
      17'd21117: data = 8'hfe;
      17'd21118: data = 8'hfe;
      17'd21119: data = 8'hfe;
      17'd21120: data = 8'h0c;
      17'd21121: data = 8'h1e;
      17'd21122: data = 8'h29;
      17'd21123: data = 8'h2d;
      17'd21124: data = 8'h39;
      17'd21125: data = 8'h40;
      17'd21126: data = 8'h3c;
      17'd21127: data = 8'h4a;
      17'd21128: data = 8'h5c;
      17'd21129: data = 8'h5f;
      17'd21130: data = 8'h64;
      17'd21131: data = 8'h6a;
      17'd21132: data = 8'h6d;
      17'd21133: data = 8'h65;
      17'd21134: data = 8'h63;
      17'd21135: data = 8'h63;
      17'd21136: data = 8'h5f;
      17'd21137: data = 8'h57;
      17'd21138: data = 8'h45;
      17'd21139: data = 8'h31;
      17'd21140: data = 8'h23;
      17'd21141: data = 8'h13;
      17'd21142: data = 8'h05;
      17'd21143: data = 8'h0a;
      17'd21144: data = 8'h13;
      17'd21145: data = 8'h12;
      17'd21146: data = 8'h12;
      17'd21147: data = 8'h15;
      17'd21148: data = 8'h0e;
      17'd21149: data = 8'h02;
      17'd21150: data = 8'hf6;
      17'd21151: data = 8'heb;
      17'd21152: data = 8'hdc;
      17'd21153: data = 8'hcd;
      17'd21154: data = 8'hbd;
      17'd21155: data = 8'hb4;
      17'd21156: data = 8'hae;
      17'd21157: data = 8'hac;
      17'd21158: data = 8'hb3;
      17'd21159: data = 8'hc1;
      17'd21160: data = 8'hcd;
      17'd21161: data = 8'hd3;
      17'd21162: data = 8'hd8;
      17'd21163: data = 8'hdc;
      17'd21164: data = 8'he0;
      17'd21165: data = 8'he4;
      17'd21166: data = 8'hed;
      17'd21167: data = 8'hfa;
      17'd21168: data = 8'h00;
      17'd21169: data = 8'h02;
      17'd21170: data = 8'h09;
      17'd21171: data = 8'h06;
      17'd21172: data = 8'h05;
      17'd21173: data = 8'h04;
      17'd21174: data = 8'h04;
      17'd21175: data = 8'h0d;
      17'd21176: data = 8'h15;
      17'd21177: data = 8'h1a;
      17'd21178: data = 8'h22;
      17'd21179: data = 8'h2d;
      17'd21180: data = 8'h3c;
      17'd21181: data = 8'h43;
      17'd21182: data = 8'h4e;
      17'd21183: data = 8'h53;
      17'd21184: data = 8'h56;
      17'd21185: data = 8'h4a;
      17'd21186: data = 8'h34;
      17'd21187: data = 8'h24;
      17'd21188: data = 8'h16;
      17'd21189: data = 8'h09;
      17'd21190: data = 8'h05;
      17'd21191: data = 8'h01;
      17'd21192: data = 8'hfd;
      17'd21193: data = 8'hf6;
      17'd21194: data = 8'hf5;
      17'd21195: data = 8'hf6;
      17'd21196: data = 8'hf1;
      17'd21197: data = 8'hed;
      17'd21198: data = 8'heb;
      17'd21199: data = 8'he5;
      17'd21200: data = 8'hdc;
      17'd21201: data = 8'hd2;
      17'd21202: data = 8'hc5;
      17'd21203: data = 8'hbc;
      17'd21204: data = 8'hb4;
      17'd21205: data = 8'hac;
      17'd21206: data = 8'hb0;
      17'd21207: data = 8'hb0;
      17'd21208: data = 8'hab;
      17'd21209: data = 8'hab;
      17'd21210: data = 8'hac;
      17'd21211: data = 8'hb0;
      17'd21212: data = 8'hb4;
      17'd21213: data = 8'hb9;
      17'd21214: data = 8'hc5;
      17'd21215: data = 8'hd2;
      17'd21216: data = 8'hda;
      17'd21217: data = 8'hde;
      17'd21218: data = 8'he2;
      17'd21219: data = 8'hde;
      17'd21220: data = 8'hde;
      17'd21221: data = 8'hdc;
      17'd21222: data = 8'hdc;
      17'd21223: data = 8'he0;
      17'd21224: data = 8'he3;
      17'd21225: data = 8'hed;
      17'd21226: data = 8'hf5;
      17'd21227: data = 8'hfe;
      17'd21228: data = 8'h0a;
      17'd21229: data = 8'h1c;
      17'd21230: data = 8'h24;
      17'd21231: data = 8'h2c;
      17'd21232: data = 8'h35;
      17'd21233: data = 8'h34;
      17'd21234: data = 8'h2d;
      17'd21235: data = 8'h26;
      17'd21236: data = 8'h27;
      17'd21237: data = 8'h1f;
      17'd21238: data = 8'h26;
      17'd21239: data = 8'h29;
      17'd21240: data = 8'h2b;
      17'd21241: data = 8'h2d;
      17'd21242: data = 8'h2c;
      17'd21243: data = 8'h2d;
      17'd21244: data = 8'h26;
      17'd21245: data = 8'h23;
      17'd21246: data = 8'h1c;
      17'd21247: data = 8'h1a;
      17'd21248: data = 8'h15;
      17'd21249: data = 8'h12;
      17'd21250: data = 8'h04;
      17'd21251: data = 8'hfd;
      17'd21252: data = 8'hfc;
      17'd21253: data = 8'hf5;
      17'd21254: data = 8'hf1;
      17'd21255: data = 8'hf1;
      17'd21256: data = 8'hf5;
      17'd21257: data = 8'heb;
      17'd21258: data = 8'he5;
      17'd21259: data = 8'hde;
      17'd21260: data = 8'he0;
      17'd21261: data = 8'hd8;
      17'd21262: data = 8'he4;
      17'd21263: data = 8'he3;
      17'd21264: data = 8'he7;
      17'd21265: data = 8'he5;
      17'd21266: data = 8'hf1;
      17'd21267: data = 8'hfe;
      17'd21268: data = 8'h00;
      17'd21269: data = 8'h0e;
      17'd21270: data = 8'h12;
      17'd21271: data = 8'hfd;
      17'd21272: data = 8'hfa;
      17'd21273: data = 8'heb;
      17'd21274: data = 8'hc0;
      17'd21275: data = 8'hbd;
      17'd21276: data = 8'hc0;
      17'd21277: data = 8'hc2;
      17'd21278: data = 8'hd6;
      17'd21279: data = 8'h05;
      17'd21280: data = 8'h22;
      17'd21281: data = 8'h2f;
      17'd21282: data = 8'h4e;
      17'd21283: data = 8'h65;
      17'd21284: data = 8'h5a;
      17'd21285: data = 8'h67;
      17'd21286: data = 8'h64;
      17'd21287: data = 8'h43;
      17'd21288: data = 8'h3e;
      17'd21289: data = 8'h1e;
      17'd21290: data = 8'h0a;
      17'd21291: data = 8'h0d;
      17'd21292: data = 8'h0d;
      17'd21293: data = 8'h1b;
      17'd21294: data = 8'h22;
      17'd21295: data = 8'h31;
      17'd21296: data = 8'h36;
      17'd21297: data = 8'h29;
      17'd21298: data = 8'h34;
      17'd21299: data = 8'h33;
      17'd21300: data = 8'h2d;
      17'd21301: data = 8'h34;
      17'd21302: data = 8'h2b;
      17'd21303: data = 8'h26;
      17'd21304: data = 8'h1a;
      17'd21305: data = 8'h01;
      17'd21306: data = 8'hef;
      17'd21307: data = 8'hdb;
      17'd21308: data = 8'hd8;
      17'd21309: data = 8'hce;
      17'd21310: data = 8'hb3;
      17'd21311: data = 8'hbb;
      17'd21312: data = 8'hae;
      17'd21313: data = 8'h9a;
      17'd21314: data = 8'ha8;
      17'd21315: data = 8'hbb;
      17'd21316: data = 8'hc2;
      17'd21317: data = 8'hce;
      17'd21318: data = 8'he0;
      17'd21319: data = 8'he0;
      17'd21320: data = 8'hd3;
      17'd21321: data = 8'hc2;
      17'd21322: data = 8'hb9;
      17'd21323: data = 8'hae;
      17'd21324: data = 8'ha6;
      17'd21325: data = 8'h9d;
      17'd21326: data = 8'h9d;
      17'd21327: data = 8'ha3;
      17'd21328: data = 8'h9d;
      17'd21329: data = 8'ha8;
      17'd21330: data = 8'hc4;
      17'd21331: data = 8'hda;
      17'd21332: data = 8'hf4;
      17'd21333: data = 8'h09;
      17'd21334: data = 8'h13;
      17'd21335: data = 8'h1e;
      17'd21336: data = 8'h22;
      17'd21337: data = 8'h24;
      17'd21338: data = 8'h2c;
      17'd21339: data = 8'h34;
      17'd21340: data = 8'h39;
      17'd21341: data = 8'h39;
      17'd21342: data = 8'h3a;
      17'd21343: data = 8'h39;
      17'd21344: data = 8'h2f;
      17'd21345: data = 8'h2f;
      17'd21346: data = 8'h34;
      17'd21347: data = 8'h39;
      17'd21348: data = 8'h40;
      17'd21349: data = 8'h46;
      17'd21350: data = 8'h52;
      17'd21351: data = 8'h52;
      17'd21352: data = 8'h53;
      17'd21353: data = 8'h5f;
      17'd21354: data = 8'h5d;
      17'd21355: data = 8'h5c;
      17'd21356: data = 8'h5b;
      17'd21357: data = 8'h47;
      17'd21358: data = 8'h34;
      17'd21359: data = 8'h22;
      17'd21360: data = 8'h04;
      17'd21361: data = 8'hf2;
      17'd21362: data = 8'he9;
      17'd21363: data = 8'he3;
      17'd21364: data = 8'hde;
      17'd21365: data = 8'he4;
      17'd21366: data = 8'hed;
      17'd21367: data = 8'heb;
      17'd21368: data = 8'hed;
      17'd21369: data = 8'hf1;
      17'd21370: data = 8'hec;
      17'd21371: data = 8'hed;
      17'd21372: data = 8'he9;
      17'd21373: data = 8'hde;
      17'd21374: data = 8'hd8;
      17'd21375: data = 8'hcd;
      17'd21376: data = 8'hc1;
      17'd21377: data = 8'hc1;
      17'd21378: data = 8'hc5;
      17'd21379: data = 8'hc6;
      17'd21380: data = 8'hc9;
      17'd21381: data = 8'hd2;
      17'd21382: data = 8'hdc;
      17'd21383: data = 8'hdc;
      17'd21384: data = 8'he4;
      17'd21385: data = 8'hf5;
      17'd21386: data = 8'h04;
      17'd21387: data = 8'h11;
      17'd21388: data = 8'h1c;
      17'd21389: data = 8'h26;
      17'd21390: data = 8'h2c;
      17'd21391: data = 8'h33;
      17'd21392: data = 8'h33;
      17'd21393: data = 8'h31;
      17'd21394: data = 8'h31;
      17'd21395: data = 8'h2b;
      17'd21396: data = 8'h22;
      17'd21397: data = 8'h23;
      17'd21398: data = 8'h1e;
      17'd21399: data = 8'h1c;
      17'd21400: data = 8'h23;
      17'd21401: data = 8'h27;
      17'd21402: data = 8'h31;
      17'd21403: data = 8'h3a;
      17'd21404: data = 8'h3e;
      17'd21405: data = 8'h39;
      17'd21406: data = 8'h34;
      17'd21407: data = 8'h29;
      17'd21408: data = 8'h1b;
      17'd21409: data = 8'h12;
      17'd21410: data = 8'h02;
      17'd21411: data = 8'hf4;
      17'd21412: data = 8'he4;
      17'd21413: data = 8'hdb;
      17'd21414: data = 8'hd2;
      17'd21415: data = 8'hcb;
      17'd21416: data = 8'hcd;
      17'd21417: data = 8'hcd;
      17'd21418: data = 8'hca;
      17'd21419: data = 8'hc9;
      17'd21420: data = 8'hca;
      17'd21421: data = 8'hc6;
      17'd21422: data = 8'hc1;
      17'd21423: data = 8'hc0;
      17'd21424: data = 8'hc4;
      17'd21425: data = 8'hc5;
      17'd21426: data = 8'hc5;
      17'd21427: data = 8'hc4;
      17'd21428: data = 8'hc1;
      17'd21429: data = 8'hc0;
      17'd21430: data = 8'hbd;
      17'd21431: data = 8'hbc;
      17'd21432: data = 8'hc2;
      17'd21433: data = 8'hc6;
      17'd21434: data = 8'hca;
      17'd21435: data = 8'hd1;
      17'd21436: data = 8'hda;
      17'd21437: data = 8'he2;
      17'd21438: data = 8'heb;
      17'd21439: data = 8'hf6;
      17'd21440: data = 8'hfd;
      17'd21441: data = 8'h04;
      17'd21442: data = 8'h09;
      17'd21443: data = 8'h0a;
      17'd21444: data = 8'h0e;
      17'd21445: data = 8'h12;
      17'd21446: data = 8'h0c;
      17'd21447: data = 8'h0d;
      17'd21448: data = 8'h16;
      17'd21449: data = 8'h16;
      17'd21450: data = 8'h1c;
      17'd21451: data = 8'h23;
      17'd21452: data = 8'h24;
      17'd21453: data = 8'h24;
      17'd21454: data = 8'h27;
      17'd21455: data = 8'h24;
      17'd21456: data = 8'h23;
      17'd21457: data = 8'h23;
      17'd21458: data = 8'h22;
      17'd21459: data = 8'h23;
      17'd21460: data = 8'h26;
      17'd21461: data = 8'h1e;
      17'd21462: data = 8'h1b;
      17'd21463: data = 8'h1e;
      17'd21464: data = 8'h12;
      17'd21465: data = 8'h12;
      17'd21466: data = 8'h0d;
      17'd21467: data = 8'h04;
      17'd21468: data = 8'h02;
      17'd21469: data = 8'hfc;
      17'd21470: data = 8'hf6;
      17'd21471: data = 8'hf4;
      17'd21472: data = 8'hf2;
      17'd21473: data = 8'hf2;
      17'd21474: data = 8'hfc;
      17'd21475: data = 8'hf6;
      17'd21476: data = 8'hf5;
      17'd21477: data = 8'hed;
      17'd21478: data = 8'hed;
      17'd21479: data = 8'he7;
      17'd21480: data = 8'he7;
      17'd21481: data = 8'hf1;
      17'd21482: data = 8'he4;
      17'd21483: data = 8'hed;
      17'd21484: data = 8'hf5;
      17'd21485: data = 8'hf5;
      17'd21486: data = 8'h02;
      17'd21487: data = 8'h13;
      17'd21488: data = 8'h16;
      17'd21489: data = 8'h1b;
      17'd21490: data = 8'h15;
      17'd21491: data = 8'h0c;
      17'd21492: data = 8'hf2;
      17'd21493: data = 8'hdb;
      17'd21494: data = 8'hc9;
      17'd21495: data = 8'hc1;
      17'd21496: data = 8'hca;
      17'd21497: data = 8'hde;
      17'd21498: data = 8'h01;
      17'd21499: data = 8'h1f;
      17'd21500: data = 8'h31;
      17'd21501: data = 8'h4b;
      17'd21502: data = 8'h5d;
      17'd21503: data = 8'h5b;
      17'd21504: data = 8'h5f;
      17'd21505: data = 8'h5a;
      17'd21506: data = 8'h4d;
      17'd21507: data = 8'h34;
      17'd21508: data = 8'h1f;
      17'd21509: data = 8'h15;
      17'd21510: data = 8'h09;
      17'd21511: data = 8'h0c;
      17'd21512: data = 8'h0d;
      17'd21513: data = 8'h15;
      17'd21514: data = 8'h1f;
      17'd21515: data = 8'h22;
      17'd21516: data = 8'h22;
      17'd21517: data = 8'h23;
      17'd21518: data = 8'h15;
      17'd21519: data = 8'h1b;
      17'd21520: data = 8'h1f;
      17'd21521: data = 8'h22;
      17'd21522: data = 8'h1c;
      17'd21523: data = 8'h15;
      17'd21524: data = 8'h12;
      17'd21525: data = 8'h04;
      17'd21526: data = 8'hfc;
      17'd21527: data = 8'hed;
      17'd21528: data = 8'hdc;
      17'd21529: data = 8'hce;
      17'd21530: data = 8'hc0;
      17'd21531: data = 8'hac;
      17'd21532: data = 8'ha4;
      17'd21533: data = 8'ha2;
      17'd21534: data = 8'haa;
      17'd21535: data = 8'hb4;
      17'd21536: data = 8'hc2;
      17'd21537: data = 8'hd8;
      17'd21538: data = 8'he5;
      17'd21539: data = 8'he4;
      17'd21540: data = 8'he4;
      17'd21541: data = 8'he3;
      17'd21542: data = 8'hd5;
      17'd21543: data = 8'hc5;
      17'd21544: data = 8'hbb;
      17'd21545: data = 8'hb3;
      17'd21546: data = 8'hab;
      17'd21547: data = 8'ha8;
      17'd21548: data = 8'hac;
      17'd21549: data = 8'hb9;
      17'd21550: data = 8'hcb;
      17'd21551: data = 8'hdc;
      17'd21552: data = 8'hf1;
      17'd21553: data = 8'h04;
      17'd21554: data = 8'h0a;
      17'd21555: data = 8'h15;
      17'd21556: data = 8'h1e;
      17'd21557: data = 8'h24;
      17'd21558: data = 8'h2c;
      17'd21559: data = 8'h34;
      17'd21560: data = 8'h3e;
      17'd21561: data = 8'h45;
      17'd21562: data = 8'h43;
      17'd21563: data = 8'h3c;
      17'd21564: data = 8'h3c;
      17'd21565: data = 8'h34;
      17'd21566: data = 8'h2d;
      17'd21567: data = 8'h2b;
      17'd21568: data = 8'h2c;
      17'd21569: data = 8'h2f;
      17'd21570: data = 8'h31;
      17'd21571: data = 8'h36;
      17'd21572: data = 8'h3e;
      17'd21573: data = 8'h47;
      17'd21574: data = 8'h4e;
      17'd21575: data = 8'h53;
      17'd21576: data = 8'h52;
      17'd21577: data = 8'h4b;
      17'd21578: data = 8'h3a;
      17'd21579: data = 8'h26;
      17'd21580: data = 8'h0e;
      17'd21581: data = 8'hfa;
      17'd21582: data = 8'hec;
      17'd21583: data = 8'he2;
      17'd21584: data = 8'hda;
      17'd21585: data = 8'hd6;
      17'd21586: data = 8'hd5;
      17'd21587: data = 8'hd8;
      17'd21588: data = 8'he0;
      17'd21589: data = 8'he3;
      17'd21590: data = 8'he4;
      17'd21591: data = 8'he7;
      17'd21592: data = 8'he7;
      17'd21593: data = 8'he4;
      17'd21594: data = 8'he0;
      17'd21595: data = 8'he0;
      17'd21596: data = 8'hde;
      17'd21597: data = 8'hde;
      17'd21598: data = 8'hdb;
      17'd21599: data = 8'hdc;
      17'd21600: data = 8'he0;
      17'd21601: data = 8'hdc;
      17'd21602: data = 8'hdc;
      17'd21603: data = 8'he4;
      17'd21604: data = 8'he9;
      17'd21605: data = 8'he9;
      17'd21606: data = 8'hf2;
      17'd21607: data = 8'hfd;
      17'd21608: data = 8'h0c;
      17'd21609: data = 8'h1a;
      17'd21610: data = 8'h27;
      17'd21611: data = 8'h36;
      17'd21612: data = 8'h3d;
      17'd21613: data = 8'h40;
      17'd21614: data = 8'h40;
      17'd21615: data = 8'h3a;
      17'd21616: data = 8'h34;
      17'd21617: data = 8'h26;
      17'd21618: data = 8'h1a;
      17'd21619: data = 8'h12;
      17'd21620: data = 8'h0a;
      17'd21621: data = 8'h09;
      17'd21622: data = 8'h0e;
      17'd21623: data = 8'h15;
      17'd21624: data = 8'h1b;
      17'd21625: data = 8'h22;
      17'd21626: data = 8'h26;
      17'd21627: data = 8'h22;
      17'd21628: data = 8'h1b;
      17'd21629: data = 8'h16;
      17'd21630: data = 8'h06;
      17'd21631: data = 8'hfd;
      17'd21632: data = 8'hf1;
      17'd21633: data = 8'he2;
      17'd21634: data = 8'hdb;
      17'd21635: data = 8'hd5;
      17'd21636: data = 8'hca;
      17'd21637: data = 8'hca;
      17'd21638: data = 8'hca;
      17'd21639: data = 8'hc6;
      17'd21640: data = 8'hc4;
      17'd21641: data = 8'hbc;
      17'd21642: data = 8'hc0;
      17'd21643: data = 8'hbd;
      17'd21644: data = 8'hc0;
      17'd21645: data = 8'hc5;
      17'd21646: data = 8'hcd;
      17'd21647: data = 8'hd5;
      17'd21648: data = 8'hdb;
      17'd21649: data = 8'he2;
      17'd21650: data = 8'he3;
      17'd21651: data = 8'hde;
      17'd21652: data = 8'hdb;
      17'd21653: data = 8'hda;
      17'd21654: data = 8'hd8;
      17'd21655: data = 8'hd6;
      17'd21656: data = 8'hd5;
      17'd21657: data = 8'hda;
      17'd21658: data = 8'he5;
      17'd21659: data = 8'hec;
      17'd21660: data = 8'hf4;
      17'd21661: data = 8'h01;
      17'd21662: data = 8'h0c;
      17'd21663: data = 8'h19;
      17'd21664: data = 8'h1b;
      17'd21665: data = 8'h1e;
      17'd21666: data = 8'h23;
      17'd21667: data = 8'h1c;
      17'd21668: data = 8'h16;
      17'd21669: data = 8'h15;
      17'd21670: data = 8'h19;
      17'd21671: data = 8'h16;
      17'd21672: data = 8'h16;
      17'd21673: data = 8'h1a;
      17'd21674: data = 8'h1a;
      17'd21675: data = 8'h15;
      17'd21676: data = 8'h19;
      17'd21677: data = 8'h19;
      17'd21678: data = 8'h15;
      17'd21679: data = 8'h15;
      17'd21680: data = 8'h13;
      17'd21681: data = 8'h15;
      17'd21682: data = 8'h1a;
      17'd21683: data = 8'h15;
      17'd21684: data = 8'h15;
      17'd21685: data = 8'h16;
      17'd21686: data = 8'h0c;
      17'd21687: data = 8'h0d;
      17'd21688: data = 8'h05;
      17'd21689: data = 8'h00;
      17'd21690: data = 8'hfa;
      17'd21691: data = 8'hf1;
      17'd21692: data = 8'heb;
      17'd21693: data = 8'he7;
      17'd21694: data = 8'hec;
      17'd21695: data = 8'hed;
      17'd21696: data = 8'heb;
      17'd21697: data = 8'hf4;
      17'd21698: data = 8'hf4;
      17'd21699: data = 8'hf4;
      17'd21700: data = 8'hfc;
      17'd21701: data = 8'h00;
      17'd21702: data = 8'hf6;
      17'd21703: data = 8'h00;
      17'd21704: data = 8'h0c;
      17'd21705: data = 8'h09;
      17'd21706: data = 8'h1b;
      17'd21707: data = 8'h1a;
      17'd21708: data = 8'h0e;
      17'd21709: data = 8'h12;
      17'd21710: data = 8'h04;
      17'd21711: data = 8'he4;
      17'd21712: data = 8'hdb;
      17'd21713: data = 8'hd3;
      17'd21714: data = 8'hc1;
      17'd21715: data = 8'hd2;
      17'd21716: data = 8'hef;
      17'd21717: data = 8'hfa;
      17'd21718: data = 8'h13;
      17'd21719: data = 8'h3a;
      17'd21720: data = 8'h46;
      17'd21721: data = 8'h53;
      17'd21722: data = 8'h60;
      17'd21723: data = 8'h56;
      17'd21724: data = 8'h52;
      17'd21725: data = 8'h40;
      17'd21726: data = 8'h23;
      17'd21727: data = 8'h15;
      17'd21728: data = 8'h0c;
      17'd21729: data = 8'hfa;
      17'd21730: data = 8'hf6;
      17'd21731: data = 8'h00;
      17'd21732: data = 8'h02;
      17'd21733: data = 8'h0a;
      17'd21734: data = 8'h12;
      17'd21735: data = 8'h1a;
      17'd21736: data = 8'h1f;
      17'd21737: data = 8'h1f;
      17'd21738: data = 8'h1c;
      17'd21739: data = 8'h1b;
      17'd21740: data = 8'h15;
      17'd21741: data = 8'h0d;
      17'd21742: data = 8'h09;
      17'd21743: data = 8'h09;
      17'd21744: data = 8'h04;
      17'd21745: data = 8'hfa;
      17'd21746: data = 8'hec;
      17'd21747: data = 8'hdc;
      17'd21748: data = 8'hd1;
      17'd21749: data = 8'hb8;
      17'd21750: data = 8'ha6;
      17'd21751: data = 8'hb1;
      17'd21752: data = 8'hab;
      17'd21753: data = 8'haa;
      17'd21754: data = 8'hbd;
      17'd21755: data = 8'hc9;
      17'd21756: data = 8'hd8;
      17'd21757: data = 8'he0;
      17'd21758: data = 8'he5;
      17'd21759: data = 8'he7;
      17'd21760: data = 8'hec;
      17'd21761: data = 8'he3;
      17'd21762: data = 8'hce;
      17'd21763: data = 8'hcb;
      17'd21764: data = 8'hb9;
      17'd21765: data = 8'ha4;
      17'd21766: data = 8'ha8;
      17'd21767: data = 8'hb0;
      17'd21768: data = 8'hb4;
      17'd21769: data = 8'hc9;
      17'd21770: data = 8'he0;
      17'd21771: data = 8'hf1;
      17'd21772: data = 8'hfd;
      17'd21773: data = 8'h05;
      17'd21774: data = 8'h13;
      17'd21775: data = 8'h1f;
      17'd21776: data = 8'h24;
      17'd21777: data = 8'h2b;
      17'd21778: data = 8'h36;
      17'd21779: data = 8'h39;
      17'd21780: data = 8'h35;
      17'd21781: data = 8'h39;
      17'd21782: data = 8'h3c;
      17'd21783: data = 8'h36;
      17'd21784: data = 8'h31;
      17'd21785: data = 8'h2d;
      17'd21786: data = 8'h2f;
      17'd21787: data = 8'h27;
      17'd21788: data = 8'h23;
      17'd21789: data = 8'h29;
      17'd21790: data = 8'h31;
      17'd21791: data = 8'h35;
      17'd21792: data = 8'h3d;
      17'd21793: data = 8'h45;
      17'd21794: data = 8'h46;
      17'd21795: data = 8'h4b;
      17'd21796: data = 8'h43;
      17'd21797: data = 8'h39;
      17'd21798: data = 8'h2b;
      17'd21799: data = 8'h1a;
      17'd21800: data = 8'h05;
      17'd21801: data = 8'hf6;
      17'd21802: data = 8'he5;
      17'd21803: data = 8'hd6;
      17'd21804: data = 8'hd1;
      17'd21805: data = 8'hcd;
      17'd21806: data = 8'hd2;
      17'd21807: data = 8'hd8;
      17'd21808: data = 8'he0;
      17'd21809: data = 8'he3;
      17'd21810: data = 8'he3;
      17'd21811: data = 8'he3;
      17'd21812: data = 8'he3;
      17'd21813: data = 8'heb;
      17'd21814: data = 8'hec;
      17'd21815: data = 8'he9;
      17'd21816: data = 8'he7;
      17'd21817: data = 8'he5;
      17'd21818: data = 8'he2;
      17'd21819: data = 8'hdc;
      17'd21820: data = 8'hdc;
      17'd21821: data = 8'hda;
      17'd21822: data = 8'hda;
      17'd21823: data = 8'hdc;
      17'd21824: data = 8'he5;
      17'd21825: data = 8'hf1;
      17'd21826: data = 8'hfd;
      17'd21827: data = 8'h0c;
      17'd21828: data = 8'h1c;
      17'd21829: data = 8'h27;
      17'd21830: data = 8'h34;
      17'd21831: data = 8'h3d;
      17'd21832: data = 8'h40;
      17'd21833: data = 8'h40;
      17'd21834: data = 8'h36;
      17'd21835: data = 8'h2d;
      17'd21836: data = 8'h22;
      17'd21837: data = 8'h16;
      17'd21838: data = 8'h0d;
      17'd21839: data = 8'h06;
      17'd21840: data = 8'h04;
      17'd21841: data = 8'hfe;
      17'd21842: data = 8'h04;
      17'd21843: data = 8'h0a;
      17'd21844: data = 8'h0d;
      17'd21845: data = 8'h0d;
      17'd21846: data = 8'h0e;
      17'd21847: data = 8'h0d;
      17'd21848: data = 8'h0c;
      17'd21849: data = 8'h06;
      17'd21850: data = 8'hfc;
      17'd21851: data = 8'hf1;
      17'd21852: data = 8'he4;
      17'd21853: data = 8'he0;
      17'd21854: data = 8'hd6;
      17'd21855: data = 8'hce;
      17'd21856: data = 8'hc9;
      17'd21857: data = 8'hc1;
      17'd21858: data = 8'hbb;
      17'd21859: data = 8'hbd;
      17'd21860: data = 8'hc0;
      17'd21861: data = 8'hb9;
      17'd21862: data = 8'hbd;
      17'd21863: data = 8'hc5;
      17'd21864: data = 8'hc9;
      17'd21865: data = 8'hce;
      17'd21866: data = 8'hd5;
      17'd21867: data = 8'hdb;
      17'd21868: data = 8'he2;
      17'd21869: data = 8'he4;
      17'd21870: data = 8'he7;
      17'd21871: data = 8'he9;
      17'd21872: data = 8'he3;
      17'd21873: data = 8'hdc;
      17'd21874: data = 8'hdb;
      17'd21875: data = 8'hda;
      17'd21876: data = 8'hdb;
      17'd21877: data = 8'he4;
      17'd21878: data = 8'he9;
      17'd21879: data = 8'hef;
      17'd21880: data = 8'hfd;
      17'd21881: data = 8'h0a;
      17'd21882: data = 8'h16;
      17'd21883: data = 8'h1c;
      17'd21884: data = 8'h22;
      17'd21885: data = 8'h24;
      17'd21886: data = 8'h26;
      17'd21887: data = 8'h23;
      17'd21888: data = 8'h1f;
      17'd21889: data = 8'h24;
      17'd21890: data = 8'h1c;
      17'd21891: data = 8'h19;
      17'd21892: data = 8'h1b;
      17'd21893: data = 8'h1b;
      17'd21894: data = 8'h19;
      17'd21895: data = 8'h19;
      17'd21896: data = 8'h15;
      17'd21897: data = 8'h11;
      17'd21898: data = 8'h11;
      17'd21899: data = 8'h0e;
      17'd21900: data = 8'h0d;
      17'd21901: data = 8'h11;
      17'd21902: data = 8'h0e;
      17'd21903: data = 8'h0e;
      17'd21904: data = 8'h11;
      17'd21905: data = 8'h0c;
      17'd21906: data = 8'h0a;
      17'd21907: data = 8'h0d;
      17'd21908: data = 8'h06;
      17'd21909: data = 8'hfe;
      17'd21910: data = 8'hfc;
      17'd21911: data = 8'hfa;
      17'd21912: data = 8'hed;
      17'd21913: data = 8'hec;
      17'd21914: data = 8'hf1;
      17'd21915: data = 8'he5;
      17'd21916: data = 8'he4;
      17'd21917: data = 8'hef;
      17'd21918: data = 8'hef;
      17'd21919: data = 8'hf2;
      17'd21920: data = 8'hfa;
      17'd21921: data = 8'hfe;
      17'd21922: data = 8'h06;
      17'd21923: data = 8'h0e;
      17'd21924: data = 8'h19;
      17'd21925: data = 8'h23;
      17'd21926: data = 8'h24;
      17'd21927: data = 8'h29;
      17'd21928: data = 8'h1c;
      17'd21929: data = 8'h1c;
      17'd21930: data = 8'h0a;
      17'd21931: data = 8'he5;
      17'd21932: data = 8'he7;
      17'd21933: data = 8'hd1;
      17'd21934: data = 8'hc4;
      17'd21935: data = 8'hd6;
      17'd21936: data = 8'he5;
      17'd21937: data = 8'hf9;
      17'd21938: data = 8'h12;
      17'd21939: data = 8'h33;
      17'd21940: data = 8'h4a;
      17'd21941: data = 8'h53;
      17'd21942: data = 8'h5d;
      17'd21943: data = 8'h5a;
      17'd21944: data = 8'h4e;
      17'd21945: data = 8'h45;
      17'd21946: data = 8'h26;
      17'd21947: data = 8'h1a;
      17'd21948: data = 8'h0d;
      17'd21949: data = 8'hf6;
      17'd21950: data = 8'hf6;
      17'd21951: data = 8'hf4;
      17'd21952: data = 8'hf2;
      17'd21953: data = 8'h02;
      17'd21954: data = 8'h06;
      17'd21955: data = 8'h12;
      17'd21956: data = 8'h16;
      17'd21957: data = 8'h1a;
      17'd21958: data = 8'h1f;
      17'd21959: data = 8'h19;
      17'd21960: data = 8'h1b;
      17'd21961: data = 8'h16;
      17'd21962: data = 8'h0c;
      17'd21963: data = 8'h0a;
      17'd21964: data = 8'h05;
      17'd21965: data = 8'h01;
      17'd21966: data = 8'hf2;
      17'd21967: data = 8'hde;
      17'd21968: data = 8'hdb;
      17'd21969: data = 8'hbd;
      17'd21970: data = 8'hb1;
      17'd21971: data = 8'hb5;
      17'd21972: data = 8'hae;
      17'd21973: data = 8'hb3;
      17'd21974: data = 8'hb8;
      17'd21975: data = 8'hc1;
      17'd21976: data = 8'hd2;
      17'd21977: data = 8'hde;
      17'd21978: data = 8'he3;
      17'd21979: data = 8'hf1;
      17'd21980: data = 8'hf5;
      17'd21981: data = 8'he9;
      17'd21982: data = 8'he2;
      17'd21983: data = 8'hdc;
      17'd21984: data = 8'hcb;
      17'd21985: data = 8'hb9;
      17'd21986: data = 8'hb5;
      17'd21987: data = 8'hb5;
      17'd21988: data = 8'hb3;
      17'd21989: data = 8'hc0;
      17'd21990: data = 8'hcd;
      17'd21991: data = 8'hde;
      17'd21992: data = 8'hf1;
      17'd21993: data = 8'hfa;
      17'd21994: data = 8'h11;
      17'd21995: data = 8'h23;
      17'd21996: data = 8'h27;
      17'd21997: data = 8'h2f;
      17'd21998: data = 8'h3c;
      17'd21999: data = 8'h3c;
      17'd22000: data = 8'h39;
      17'd22001: data = 8'h3c;
      17'd22002: data = 8'h40;
      17'd22003: data = 8'h39;
      17'd22004: data = 8'h31;
      17'd22005: data = 8'h31;
      17'd22006: data = 8'h27;
      17'd22007: data = 8'h23;
      17'd22008: data = 8'h22;
      17'd22009: data = 8'h23;
      17'd22010: data = 8'h29;
      17'd22011: data = 8'h2c;
      17'd22012: data = 8'h34;
      17'd22013: data = 8'h3c;
      17'd22014: data = 8'h3d;
      17'd22015: data = 8'h42;
      17'd22016: data = 8'h40;
      17'd22017: data = 8'h3c;
      17'd22018: data = 8'h35;
      17'd22019: data = 8'h26;
      17'd22020: data = 8'h19;
      17'd22021: data = 8'h06;
      17'd22022: data = 8'hf5;
      17'd22023: data = 8'he5;
      17'd22024: data = 8'hd6;
      17'd22025: data = 8'hd1;
      17'd22026: data = 8'hd1;
      17'd22027: data = 8'hce;
      17'd22028: data = 8'hd2;
      17'd22029: data = 8'hd8;
      17'd22030: data = 8'he0;
      17'd22031: data = 8'he4;
      17'd22032: data = 8'heb;
      17'd22033: data = 8'hf2;
      17'd22034: data = 8'hf2;
      17'd22035: data = 8'hed;
      17'd22036: data = 8'hed;
      17'd22037: data = 8'hed;
      17'd22038: data = 8'he9;
      17'd22039: data = 8'he4;
      17'd22040: data = 8'he3;
      17'd22041: data = 8'he2;
      17'd22042: data = 8'hdc;
      17'd22043: data = 8'hdc;
      17'd22044: data = 8'he3;
      17'd22045: data = 8'he9;
      17'd22046: data = 8'hed;
      17'd22047: data = 8'hf6;
      17'd22048: data = 8'h04;
      17'd22049: data = 8'h12;
      17'd22050: data = 8'h1a;
      17'd22051: data = 8'h26;
      17'd22052: data = 8'h33;
      17'd22053: data = 8'h35;
      17'd22054: data = 8'h39;
      17'd22055: data = 8'h36;
      17'd22056: data = 8'h31;
      17'd22057: data = 8'h29;
      17'd22058: data = 8'h1c;
      17'd22059: data = 8'h12;
      17'd22060: data = 8'h09;
      17'd22061: data = 8'hfe;
      17'd22062: data = 8'hf9;
      17'd22063: data = 8'hf5;
      17'd22064: data = 8'hf5;
      17'd22065: data = 8'hf9;
      17'd22066: data = 8'h01;
      17'd22067: data = 8'h0c;
      17'd22068: data = 8'h06;
      17'd22069: data = 8'h05;
      17'd22070: data = 8'h05;
      17'd22071: data = 8'h00;
      17'd22072: data = 8'hfa;
      17'd22073: data = 8'hef;
      17'd22074: data = 8'he3;
      17'd22075: data = 8'hd6;
      17'd22076: data = 8'hce;
      17'd22077: data = 8'hc6;
      17'd22078: data = 8'hc1;
      17'd22079: data = 8'hc0;
      17'd22080: data = 8'hbd;
      17'd22081: data = 8'hbc;
      17'd22082: data = 8'hbc;
      17'd22083: data = 8'hc1;
      17'd22084: data = 8'hc5;
      17'd22085: data = 8'hcb;
      17'd22086: data = 8'hd1;
      17'd22087: data = 8'hd8;
      17'd22088: data = 8'hdc;
      17'd22089: data = 8'he0;
      17'd22090: data = 8'he9;
      17'd22091: data = 8'hec;
      17'd22092: data = 8'hed;
      17'd22093: data = 8'hec;
      17'd22094: data = 8'he7;
      17'd22095: data = 8'he3;
      17'd22096: data = 8'he3;
      17'd22097: data = 8'he2;
      17'd22098: data = 8'he2;
      17'd22099: data = 8'he7;
      17'd22100: data = 8'hed;
      17'd22101: data = 8'hf6;
      17'd22102: data = 8'h04;
      17'd22103: data = 8'h11;
      17'd22104: data = 8'h16;
      17'd22105: data = 8'h1e;
      17'd22106: data = 8'h23;
      17'd22107: data = 8'h2b;
      17'd22108: data = 8'h29;
      17'd22109: data = 8'h29;
      17'd22110: data = 8'h27;
      17'd22111: data = 8'h23;
      17'd22112: data = 8'h1f;
      17'd22113: data = 8'h1a;
      17'd22114: data = 8'h16;
      17'd22115: data = 8'h12;
      17'd22116: data = 8'h11;
      17'd22117: data = 8'h0d;
      17'd22118: data = 8'h0a;
      17'd22119: data = 8'h0e;
      17'd22120: data = 8'h0a;
      17'd22121: data = 8'h12;
      17'd22122: data = 8'h0e;
      17'd22123: data = 8'h0c;
      17'd22124: data = 8'h13;
      17'd22125: data = 8'h12;
      17'd22126: data = 8'h0d;
      17'd22127: data = 8'h15;
      17'd22128: data = 8'h13;
      17'd22129: data = 8'h0a;
      17'd22130: data = 8'h11;
      17'd22131: data = 8'h06;
      17'd22132: data = 8'hfe;
      17'd22133: data = 8'hfd;
      17'd22134: data = 8'hf5;
      17'd22135: data = 8'he7;
      17'd22136: data = 8'hec;
      17'd22137: data = 8'he7;
      17'd22138: data = 8'he4;
      17'd22139: data = 8'hf1;
      17'd22140: data = 8'hf5;
      17'd22141: data = 8'hf5;
      17'd22142: data = 8'h06;
      17'd22143: data = 8'h0e;
      17'd22144: data = 8'h11;
      17'd22145: data = 8'h27;
      17'd22146: data = 8'h2c;
      17'd22147: data = 8'h2b;
      17'd22148: data = 8'h2c;
      17'd22149: data = 8'h1c;
      17'd22150: data = 8'h09;
      17'd22151: data = 8'hfe;
      17'd22152: data = 8'he0;
      17'd22153: data = 8'hce;
      17'd22154: data = 8'hd1;
      17'd22155: data = 8'hc9;
      17'd22156: data = 8'hce;
      17'd22157: data = 8'hf1;
      17'd22158: data = 8'hfe;
      17'd22159: data = 8'h0e;
      17'd22160: data = 8'h2f;
      17'd22161: data = 8'h3e;
      17'd22162: data = 8'h4b;
      17'd22163: data = 8'h56;
      17'd22164: data = 8'h52;
      17'd22165: data = 8'h45;
      17'd22166: data = 8'h42;
      17'd22167: data = 8'h27;
      17'd22168: data = 8'h16;
      17'd22169: data = 8'h11;
      17'd22170: data = 8'h00;
      17'd22171: data = 8'hf4;
      17'd22172: data = 8'hf9;
      17'd22173: data = 8'hfa;
      17'd22174: data = 8'hf9;
      17'd22175: data = 8'h02;
      17'd22176: data = 8'h06;
      17'd22177: data = 8'h0e;
      17'd22178: data = 8'h19;
      17'd22179: data = 8'h16;
      17'd22180: data = 8'h1a;
      17'd22181: data = 8'h1e;
      17'd22182: data = 8'h13;
      17'd22183: data = 8'h12;
      17'd22184: data = 8'h12;
      17'd22185: data = 8'h0a;
      17'd22186: data = 8'h04;
      17'd22187: data = 8'hf9;
      17'd22188: data = 8'he7;
      17'd22189: data = 8'hde;
      17'd22190: data = 8'hc6;
      17'd22191: data = 8'hb4;
      17'd22192: data = 8'hb4;
      17'd22193: data = 8'hae;
      17'd22194: data = 8'haa;
      17'd22195: data = 8'hb3;
      17'd22196: data = 8'hc1;
      17'd22197: data = 8'hc6;
      17'd22198: data = 8'hd5;
      17'd22199: data = 8'he3;
      17'd22200: data = 8'heb;
      17'd22201: data = 8'hed;
      17'd22202: data = 8'hec;
      17'd22203: data = 8'he5;
      17'd22204: data = 8'he3;
      17'd22205: data = 8'hd2;
      17'd22206: data = 8'hc2;
      17'd22207: data = 8'hc4;
      17'd22208: data = 8'hbc;
      17'd22209: data = 8'hb4;
      17'd22210: data = 8'hbd;
      17'd22211: data = 8'hc9;
      17'd22212: data = 8'hd5;
      17'd22213: data = 8'he7;
      17'd22214: data = 8'hfa;
      17'd22215: data = 8'h0d;
      17'd22216: data = 8'h1f;
      17'd22217: data = 8'h27;
      17'd22218: data = 8'h33;
      17'd22219: data = 8'h43;
      17'd22220: data = 8'h40;
      17'd22221: data = 8'h40;
      17'd22222: data = 8'h45;
      17'd22223: data = 8'h43;
      17'd22224: data = 8'h3c;
      17'd22225: data = 8'h39;
      17'd22226: data = 8'h35;
      17'd22227: data = 8'h2c;
      17'd22228: data = 8'h23;
      17'd22229: data = 8'h1f;
      17'd22230: data = 8'h1f;
      17'd22231: data = 8'h22;
      17'd22232: data = 8'h22;
      17'd22233: data = 8'h27;
      17'd22234: data = 8'h33;
      17'd22235: data = 8'h33;
      17'd22236: data = 8'h35;
      17'd22237: data = 8'h39;
      17'd22238: data = 8'h3a;
      17'd22239: data = 8'h35;
      17'd22240: data = 8'h2c;
      17'd22241: data = 8'h1f;
      17'd22242: data = 8'h12;
      17'd22243: data = 8'h02;
      17'd22244: data = 8'hf1;
      17'd22245: data = 8'he3;
      17'd22246: data = 8'hd6;
      17'd22247: data = 8'hcb;
      17'd22248: data = 8'hcb;
      17'd22249: data = 8'hd1;
      17'd22250: data = 8'hd1;
      17'd22251: data = 8'hda;
      17'd22252: data = 8'he0;
      17'd22253: data = 8'he7;
      17'd22254: data = 8'hed;
      17'd22255: data = 8'hf1;
      17'd22256: data = 8'hf6;
      17'd22257: data = 8'hf9;
      17'd22258: data = 8'hf5;
      17'd22259: data = 8'hf4;
      17'd22260: data = 8'hf6;
      17'd22261: data = 8'hf5;
      17'd22262: data = 8'hed;
      17'd22263: data = 8'hec;
      17'd22264: data = 8'heb;
      17'd22265: data = 8'he7;
      17'd22266: data = 8'he7;
      17'd22267: data = 8'heb;
      17'd22268: data = 8'hef;
      17'd22269: data = 8'hf6;
      17'd22270: data = 8'h00;
      17'd22271: data = 8'h06;
      17'd22272: data = 8'h15;
      17'd22273: data = 8'h1e;
      17'd22274: data = 8'h26;
      17'd22275: data = 8'h31;
      17'd22276: data = 8'h35;
      17'd22277: data = 8'h35;
      17'd22278: data = 8'h33;
      17'd22279: data = 8'h2c;
      17'd22280: data = 8'h23;
      17'd22281: data = 8'h19;
      17'd22282: data = 8'h0a;
      17'd22283: data = 8'h01;
      17'd22284: data = 8'hf6;
      17'd22285: data = 8'hed;
      17'd22286: data = 8'hed;
      17'd22287: data = 8'hed;
      17'd22288: data = 8'hef;
      17'd22289: data = 8'hf2;
      17'd22290: data = 8'hf9;
      17'd22291: data = 8'hfc;
      17'd22292: data = 8'hfa;
      17'd22293: data = 8'hf9;
      17'd22294: data = 8'hf6;
      17'd22295: data = 8'hf4;
      17'd22296: data = 8'he7;
      17'd22297: data = 8'hde;
      17'd22298: data = 8'hda;
      17'd22299: data = 8'hcb;
      17'd22300: data = 8'hc5;
      17'd22301: data = 8'hc1;
      17'd22302: data = 8'hbc;
      17'd22303: data = 8'hbb;
      17'd22304: data = 8'hbb;
      17'd22305: data = 8'hc0;
      17'd22306: data = 8'hc2;
      17'd22307: data = 8'hc6;
      17'd22308: data = 8'hcd;
      17'd22309: data = 8'hd6;
      17'd22310: data = 8'he2;
      17'd22311: data = 8'he5;
      17'd22312: data = 8'hef;
      17'd22313: data = 8'hf4;
      17'd22314: data = 8'hf2;
      17'd22315: data = 8'hf4;
      17'd22316: data = 8'hf5;
      17'd22317: data = 8'hf2;
      17'd22318: data = 8'hf1;
      17'd22319: data = 8'hf2;
      17'd22320: data = 8'hed;
      17'd22321: data = 8'hed;
      17'd22322: data = 8'hf1;
      17'd22323: data = 8'hf4;
      17'd22324: data = 8'hfd;
      17'd22325: data = 8'h02;
      17'd22326: data = 8'h0d;
      17'd22327: data = 8'h16;
      17'd22328: data = 8'h1f;
      17'd22329: data = 8'h27;
      17'd22330: data = 8'h2c;
      17'd22331: data = 8'h2d;
      17'd22332: data = 8'h2c;
      17'd22333: data = 8'h2c;
      17'd22334: data = 8'h27;
      17'd22335: data = 8'h22;
      17'd22336: data = 8'h1c;
      17'd22337: data = 8'h15;
      17'd22338: data = 8'h12;
      17'd22339: data = 8'h0d;
      17'd22340: data = 8'h09;
      17'd22341: data = 8'h09;
      17'd22342: data = 8'h05;
      17'd22343: data = 8'h05;
      17'd22344: data = 8'h04;
      17'd22345: data = 8'h06;
      17'd22346: data = 8'h09;
      17'd22347: data = 8'h0a;
      17'd22348: data = 8'h0c;
      17'd22349: data = 8'h0d;
      17'd22350: data = 8'h13;
      17'd22351: data = 8'h11;
      17'd22352: data = 8'h0c;
      17'd22353: data = 8'h11;
      17'd22354: data = 8'h06;
      17'd22355: data = 8'h00;
      17'd22356: data = 8'h02;
      17'd22357: data = 8'hf9;
      17'd22358: data = 8'hef;
      17'd22359: data = 8'hef;
      17'd22360: data = 8'heb;
      17'd22361: data = 8'heb;
      17'd22362: data = 8'hf2;
      17'd22363: data = 8'hf6;
      17'd22364: data = 8'hfd;
      17'd22365: data = 8'h0c;
      17'd22366: data = 8'h12;
      17'd22367: data = 8'h1b;
      17'd22368: data = 8'h2c;
      17'd22369: data = 8'h29;
      17'd22370: data = 8'h27;
      17'd22371: data = 8'h2d;
      17'd22372: data = 8'h1c;
      17'd22373: data = 8'h0a;
      17'd22374: data = 8'h01;
      17'd22375: data = 8'heb;
      17'd22376: data = 8'hda;
      17'd22377: data = 8'hd6;
      17'd22378: data = 8'hce;
      17'd22379: data = 8'hd3;
      17'd22380: data = 8'he7;
      17'd22381: data = 8'hf6;
      17'd22382: data = 8'h0a;
      17'd22383: data = 8'h24;
      17'd22384: data = 8'h35;
      17'd22385: data = 8'h42;
      17'd22386: data = 8'h4b;
      17'd22387: data = 8'h47;
      17'd22388: data = 8'h47;
      17'd22389: data = 8'h40;
      17'd22390: data = 8'h2c;
      17'd22391: data = 8'h1f;
      17'd22392: data = 8'h1c;
      17'd22393: data = 8'h0a;
      17'd22394: data = 8'h00;
      17'd22395: data = 8'hfe;
      17'd22396: data = 8'hfa;
      17'd22397: data = 8'hfa;
      17'd22398: data = 8'hfc;
      17'd22399: data = 8'h01;
      17'd22400: data = 8'h0a;
      17'd22401: data = 8'h0a;
      17'd22402: data = 8'h0e;
      17'd22403: data = 8'h15;
      17'd22404: data = 8'h19;
      17'd22405: data = 8'h11;
      17'd22406: data = 8'h19;
      17'd22407: data = 8'h1a;
      17'd22408: data = 8'h0e;
      17'd22409: data = 8'h0c;
      17'd22410: data = 8'h04;
      17'd22411: data = 8'hfa;
      17'd22412: data = 8'he3;
      17'd22413: data = 8'hd5;
      17'd22414: data = 8'hc9;
      17'd22415: data = 8'hbb;
      17'd22416: data = 8'hb0;
      17'd22417: data = 8'hab;
      17'd22418: data = 8'hb3;
      17'd22419: data = 8'hb5;
      17'd22420: data = 8'hbd;
      17'd22421: data = 8'hcd;
      17'd22422: data = 8'hdb;
      17'd22423: data = 8'he3;
      17'd22424: data = 8'he7;
      17'd22425: data = 8'heb;
      17'd22426: data = 8'heb;
      17'd22427: data = 8'he4;
      17'd22428: data = 8'hdb;
      17'd22429: data = 8'hd6;
      17'd22430: data = 8'hd5;
      17'd22431: data = 8'hcb;
      17'd22432: data = 8'hcb;
      17'd22433: data = 8'hce;
      17'd22434: data = 8'hd2;
      17'd22435: data = 8'hdc;
      17'd22436: data = 8'he7;
      17'd22437: data = 8'hf6;
      17'd22438: data = 8'h04;
      17'd22439: data = 8'h0e;
      17'd22440: data = 8'h1b;
      17'd22441: data = 8'h29;
      17'd22442: data = 8'h2f;
      17'd22443: data = 8'h35;
      17'd22444: data = 8'h3d;
      17'd22445: data = 8'h45;
      17'd22446: data = 8'h46;
      17'd22447: data = 8'h45;
      17'd22448: data = 8'h46;
      17'd22449: data = 8'h42;
      17'd22450: data = 8'h3c;
      17'd22451: data = 8'h33;
      17'd22452: data = 8'h29;
      17'd22453: data = 8'h24;
      17'd22454: data = 8'h1b;
      17'd22455: data = 8'h16;
      17'd22456: data = 8'h19;
      17'd22457: data = 8'h1b;
      17'd22458: data = 8'h1e;
      17'd22459: data = 8'h26;
      17'd22460: data = 8'h2d;
      17'd22461: data = 8'h2d;
      17'd22462: data = 8'h2c;
      17'd22463: data = 8'h29;
      17'd22464: data = 8'h1f;
      17'd22465: data = 8'h16;
      17'd22466: data = 8'h09;
      17'd22467: data = 8'hfe;
      17'd22468: data = 8'hf5;
      17'd22469: data = 8'heb;
      17'd22470: data = 8'hdc;
      17'd22471: data = 8'hd8;
      17'd22472: data = 8'hd5;
      17'd22473: data = 8'hd2;
      17'd22474: data = 8'hd2;
      17'd22475: data = 8'hd6;
      17'd22476: data = 8'hdb;
      17'd22477: data = 8'hdb;
      17'd22478: data = 8'he2;
      17'd22479: data = 8'he5;
      17'd22480: data = 8'he9;
      17'd22481: data = 8'hec;
      17'd22482: data = 8'hf2;
      17'd22483: data = 8'hf6;
      17'd22484: data = 8'hfa;
      17'd22485: data = 8'hfd;
      17'd22486: data = 8'hfe;
      17'd22487: data = 8'hfd;
      17'd22488: data = 8'hfa;
      17'd22489: data = 8'hf5;
      17'd22490: data = 8'hf2;
      17'd22491: data = 8'hf1;
      17'd22492: data = 8'hed;
      17'd22493: data = 8'hf1;
      17'd22494: data = 8'hf6;
      17'd22495: data = 8'hfd;
      17'd22496: data = 8'h05;
      17'd22497: data = 8'h13;
      17'd22498: data = 8'h1e;
      17'd22499: data = 8'h27;
      17'd22500: data = 8'h2d;
      17'd22501: data = 8'h2f;
      17'd22502: data = 8'h2d;
      17'd22503: data = 8'h29;
      17'd22504: data = 8'h22;
      17'd22505: data = 8'h19;
      17'd22506: data = 8'h0e;
      17'd22507: data = 8'h05;
      17'd22508: data = 8'hfc;
      17'd22509: data = 8'hf5;
      17'd22510: data = 8'hf1;
      17'd22511: data = 8'hec;
      17'd22512: data = 8'hec;
      17'd22513: data = 8'hed;
      17'd22514: data = 8'hed;
      17'd22515: data = 8'hed;
      17'd22516: data = 8'hec;
      17'd22517: data = 8'he9;
      17'd22518: data = 8'he7;
      17'd22519: data = 8'he5;
      17'd22520: data = 8'he3;
      17'd22521: data = 8'he2;
      17'd22522: data = 8'he0;
      17'd22523: data = 8'hdb;
      17'd22524: data = 8'hd8;
      17'd22525: data = 8'hd3;
      17'd22526: data = 8'hce;
      17'd22527: data = 8'hcd;
      17'd22528: data = 8'hca;
      17'd22529: data = 8'hc6;
      17'd22530: data = 8'hc6;
      17'd22531: data = 8'hc9;
      17'd22532: data = 8'hcd;
      17'd22533: data = 8'hd3;
      17'd22534: data = 8'hd8;
      17'd22535: data = 8'he0;
      17'd22536: data = 8'he7;
      17'd22537: data = 8'hed;
      17'd22538: data = 8'hf1;
      17'd22539: data = 8'hf4;
      17'd22540: data = 8'hf5;
      17'd22541: data = 8'hf6;
      17'd22542: data = 8'hf5;
      17'd22543: data = 8'hfa;
      17'd22544: data = 8'hfc;
      17'd22545: data = 8'hfc;
      17'd22546: data = 8'h00;
      17'd22547: data = 8'h01;
      17'd22548: data = 8'h06;
      17'd22549: data = 8'h0c;
      17'd22550: data = 8'h0e;
      17'd22551: data = 8'h12;
      17'd22552: data = 8'h15;
      17'd22553: data = 8'h13;
      17'd22554: data = 8'h1a;
      17'd22555: data = 8'h1f;
      17'd22556: data = 8'h1f;
      17'd22557: data = 8'h1f;
      17'd22558: data = 8'h23;
      17'd22559: data = 8'h23;
      17'd22560: data = 8'h23;
      17'd22561: data = 8'h1f;
      17'd22562: data = 8'h1f;
      17'd22563: data = 8'h1a;
      17'd22564: data = 8'h12;
      17'd22565: data = 8'h11;
      17'd22566: data = 8'h05;
      17'd22567: data = 8'h04;
      17'd22568: data = 8'h02;
      17'd22569: data = 8'hfe;
      17'd22570: data = 8'h01;
      17'd22571: data = 8'h01;
      17'd22572: data = 8'h06;
      17'd22573: data = 8'h06;
      17'd22574: data = 8'h0a;
      17'd22575: data = 8'h0e;
      17'd22576: data = 8'h0a;
      17'd22577: data = 8'h0d;
      17'd22578: data = 8'h06;
      17'd22579: data = 8'h05;
      17'd22580: data = 8'h05;
      17'd22581: data = 8'hf9;
      17'd22582: data = 8'hf9;
      17'd22583: data = 8'hfc;
      17'd22584: data = 8'hf2;
      17'd22585: data = 8'hf4;
      17'd22586: data = 8'hf6;
      17'd22587: data = 8'hf9;
      17'd22588: data = 8'hfc;
      17'd22589: data = 8'h01;
      17'd22590: data = 8'h0a;
      17'd22591: data = 8'h0d;
      17'd22592: data = 8'h13;
      17'd22593: data = 8'h15;
      17'd22594: data = 8'h1e;
      17'd22595: data = 8'h1a;
      17'd22596: data = 8'h16;
      17'd22597: data = 8'h0c;
      17'd22598: data = 8'h01;
      17'd22599: data = 8'hfa;
      17'd22600: data = 8'he2;
      17'd22601: data = 8'he9;
      17'd22602: data = 8'hde;
      17'd22603: data = 8'hde;
      17'd22604: data = 8'hed;
      17'd22605: data = 8'hf2;
      17'd22606: data = 8'h02;
      17'd22607: data = 8'h0d;
      17'd22608: data = 8'h1a;
      17'd22609: data = 8'h2c;
      17'd22610: data = 8'h2d;
      17'd22611: data = 8'h33;
      17'd22612: data = 8'h35;
      17'd22613: data = 8'h34;
      17'd22614: data = 8'h31;
      17'd22615: data = 8'h29;
      17'd22616: data = 8'h27;
      17'd22617: data = 8'h24;
      17'd22618: data = 8'h1c;
      17'd22619: data = 8'h15;
      17'd22620: data = 8'h11;
      17'd22621: data = 8'h09;
      17'd22622: data = 8'h04;
      17'd22623: data = 8'hfd;
      17'd22624: data = 8'hfc;
      17'd22625: data = 8'h01;
      17'd22626: data = 8'hfa;
      17'd22627: data = 8'h00;
      17'd22628: data = 8'h05;
      17'd22629: data = 8'h0a;
      17'd22630: data = 8'h15;
      17'd22631: data = 8'h0e;
      17'd22632: data = 8'h13;
      17'd22633: data = 8'h11;
      17'd22634: data = 8'h04;
      17'd22635: data = 8'hfe;
      17'd22636: data = 8'hef;
      17'd22637: data = 8'he0;
      17'd22638: data = 8'hd2;
      17'd22639: data = 8'hca;
      17'd22640: data = 8'hc5;
      17'd22641: data = 8'hbc;
      17'd22642: data = 8'hbc;
      17'd22643: data = 8'hbd;
      17'd22644: data = 8'hbd;
      17'd22645: data = 8'hc0;
      17'd22646: data = 8'hc2;
      17'd22647: data = 8'hc4;
      17'd22648: data = 8'hc6;
      17'd22649: data = 8'hca;
      17'd22650: data = 8'hca;
      17'd22651: data = 8'hd1;
      17'd22652: data = 8'hd6;
      17'd22653: data = 8'he2;
      17'd22654: data = 8'he9;
      17'd22655: data = 8'hed;
      17'd22656: data = 8'hf1;
      17'd22657: data = 8'hf4;
      17'd22658: data = 8'hf5;
      17'd22659: data = 8'hf4;
      17'd22660: data = 8'hf9;
      17'd22661: data = 8'hf9;
      17'd22662: data = 8'hfc;
      17'd22663: data = 8'h01;
      17'd22664: data = 8'h05;
      17'd22665: data = 8'h11;
      17'd22666: data = 8'h1a;
      17'd22667: data = 8'h27;
      17'd22668: data = 8'h33;
      17'd22669: data = 8'h3d;
      17'd22670: data = 8'h46;
      17'd22671: data = 8'h4a;
      17'd22672: data = 8'h47;
      17'd22673: data = 8'h45;
      17'd22674: data = 8'h45;
      17'd22675: data = 8'h42;
      17'd22676: data = 8'h3a;
      17'd22677: data = 8'h36;
      17'd22678: data = 8'h34;
      17'd22679: data = 8'h2c;
      17'd22680: data = 8'h27;
      17'd22681: data = 8'h24;
      17'd22682: data = 8'h1b;
      17'd22683: data = 8'h15;
      17'd22684: data = 8'h11;
      17'd22685: data = 8'h09;
      17'd22686: data = 8'h05;
      17'd22687: data = 8'h02;
      17'd22688: data = 8'h02;
      17'd22689: data = 8'h02;
      17'd22690: data = 8'h01;
      17'd22691: data = 8'h02;
      17'd22692: data = 8'h01;
      17'd22693: data = 8'hfd;
      17'd22694: data = 8'hf6;
      17'd22695: data = 8'hf2;
      17'd22696: data = 8'heb;
      17'd22697: data = 8'he3;
      17'd22698: data = 8'hdb;
      17'd22699: data = 8'hd8;
      17'd22700: data = 8'hd3;
      17'd22701: data = 8'hd2;
      17'd22702: data = 8'hd3;
      17'd22703: data = 8'hd5;
      17'd22704: data = 8'hda;
      17'd22705: data = 8'hde;
      17'd22706: data = 8'he5;
      17'd22707: data = 8'heb;
      17'd22708: data = 8'hed;
      17'd22709: data = 8'hf5;
      17'd22710: data = 8'hf9;
      17'd22711: data = 8'hfd;
      17'd22712: data = 8'h00;
      17'd22713: data = 8'h04;
      17'd22714: data = 8'h06;
      17'd22715: data = 8'h09;
      17'd22716: data = 8'h0d;
      17'd22717: data = 8'h11;
      17'd22718: data = 8'h13;
      17'd22719: data = 8'h13;
      17'd22720: data = 8'h13;
      17'd22721: data = 8'h13;
      17'd22722: data = 8'h12;
      17'd22723: data = 8'h0e;
      17'd22724: data = 8'h0d;
      17'd22725: data = 8'h0e;
      17'd22726: data = 8'h0d;
      17'd22727: data = 8'h11;
      17'd22728: data = 8'h12;
      17'd22729: data = 8'h13;
      17'd22730: data = 8'h16;
      17'd22731: data = 8'h12;
      17'd22732: data = 8'h11;
      17'd22733: data = 8'h0d;
      17'd22734: data = 8'h05;
      17'd22735: data = 8'h01;
      17'd22736: data = 8'hfa;
      17'd22737: data = 8'hf2;
      17'd22738: data = 8'heb;
      17'd22739: data = 8'he4;
      17'd22740: data = 8'hdc;
      17'd22741: data = 8'hd8;
      17'd22742: data = 8'hd3;
      17'd22743: data = 8'hce;
      17'd22744: data = 8'hcd;
      17'd22745: data = 8'hce;
      17'd22746: data = 8'hce;
      17'd22747: data = 8'hd1;
      17'd22748: data = 8'hd1;
      17'd22749: data = 8'hd2;
      17'd22750: data = 8'hd5;
      17'd22751: data = 8'hd6;
      17'd22752: data = 8'hd8;
      17'd22753: data = 8'hdb;
      17'd22754: data = 8'hde;
      17'd22755: data = 8'he0;
      17'd22756: data = 8'he0;
      17'd22757: data = 8'he0;
      17'd22758: data = 8'he0;
      17'd22759: data = 8'he2;
      17'd22760: data = 8'he3;
      17'd22761: data = 8'he5;
      17'd22762: data = 8'he9;
      17'd22763: data = 8'heb;
      17'd22764: data = 8'hef;
      17'd22765: data = 8'hf2;
      17'd22766: data = 8'hf4;
      17'd22767: data = 8'hfc;
      17'd22768: data = 8'h00;
      17'd22769: data = 8'h02;
      17'd22770: data = 8'h0a;
      17'd22771: data = 8'h11;
      17'd22772: data = 8'h12;
      17'd22773: data = 8'h11;
      17'd22774: data = 8'h16;
      17'd22775: data = 8'h19;
      17'd22776: data = 8'h15;
      17'd22777: data = 8'h19;
      17'd22778: data = 8'h16;
      17'd22779: data = 8'h15;
      17'd22780: data = 8'h15;
      17'd22781: data = 8'h15;
      17'd22782: data = 8'h13;
      17'd22783: data = 8'h11;
      17'd22784: data = 8'h11;
      17'd22785: data = 8'h0d;
      17'd22786: data = 8'h0e;
      17'd22787: data = 8'h0c;
      17'd22788: data = 8'h0d;
      17'd22789: data = 8'h0d;
      17'd22790: data = 8'h0c;
      17'd22791: data = 8'h0a;
      17'd22792: data = 8'h0a;
      17'd22793: data = 8'h0c;
      17'd22794: data = 8'h06;
      17'd22795: data = 8'h0c;
      17'd22796: data = 8'h0a;
      17'd22797: data = 8'h05;
      17'd22798: data = 8'h09;
      17'd22799: data = 8'h00;
      17'd22800: data = 8'hfc;
      17'd22801: data = 8'hfa;
      17'd22802: data = 8'hfd;
      17'd22803: data = 8'hfa;
      17'd22804: data = 8'hfa;
      17'd22805: data = 8'hfd;
      17'd22806: data = 8'hfa;
      17'd22807: data = 8'hf9;
      17'd22808: data = 8'hf6;
      17'd22809: data = 8'hfa;
      17'd22810: data = 8'hf9;
      17'd22811: data = 8'hfe;
      17'd22812: data = 8'h00;
      17'd22813: data = 8'h04;
      17'd22814: data = 8'h06;
      17'd22815: data = 8'h0a;
      17'd22816: data = 8'h16;
      17'd22817: data = 8'h1c;
      17'd22818: data = 8'h1e;
      17'd22819: data = 8'h0e;
      17'd22820: data = 8'h12;
      17'd22821: data = 8'h02;
      17'd22822: data = 8'heb;
      17'd22823: data = 8'he5;
      17'd22824: data = 8'he0;
      17'd22825: data = 8'he0;
      17'd22826: data = 8'hde;
      17'd22827: data = 8'hec;
      17'd22828: data = 8'hf4;
      17'd22829: data = 8'hf9;
      17'd22830: data = 8'h01;
      17'd22831: data = 8'h0e;
      17'd22832: data = 8'h1c;
      17'd22833: data = 8'h1f;
      17'd22834: data = 8'h2d;
      17'd22835: data = 8'h35;
      17'd22836: data = 8'h39;
      17'd22837: data = 8'h36;
      17'd22838: data = 8'h33;
      17'd22839: data = 8'h3e;
      17'd22840: data = 8'h35;
      17'd22841: data = 8'h2d;
      17'd22842: data = 8'h2c;
      17'd22843: data = 8'h1f;
      17'd22844: data = 8'h0e;
      17'd22845: data = 8'hfc;
      17'd22846: data = 8'hfd;
      17'd22847: data = 8'hf9;
      17'd22848: data = 8'hf1;
      17'd22849: data = 8'hf1;
      17'd22850: data = 8'hf9;
      17'd22851: data = 8'h00;
      17'd22852: data = 8'hfd;
      17'd22853: data = 8'hfe;
      17'd22854: data = 8'h05;
      17'd22855: data = 8'h09;
      17'd22856: data = 8'hfe;
      17'd22857: data = 8'hfe;
      17'd22858: data = 8'h01;
      17'd22859: data = 8'hf4;
      17'd22860: data = 8'he9;
      17'd22861: data = 8'he2;
      17'd22862: data = 8'he2;
      17'd22863: data = 8'hd3;
      17'd22864: data = 8'hc9;
      17'd22865: data = 8'hc5;
      17'd22866: data = 8'hb8;
      17'd22867: data = 8'hac;
      17'd22868: data = 8'ha6;
      17'd22869: data = 8'hab;
      17'd22870: data = 8'hac;
      17'd22871: data = 8'hae;
      17'd22872: data = 8'hbc;
      17'd22873: data = 8'hc5;
      17'd22874: data = 8'hce;
      17'd22875: data = 8'hd6;
      17'd22876: data = 8'he5;
      17'd22877: data = 8'hf1;
      17'd22878: data = 8'hf6;
      17'd22879: data = 8'hfd;
      17'd22880: data = 8'h05;
      17'd22881: data = 8'h0a;
      17'd22882: data = 8'h0c;
      17'd22883: data = 8'h12;
      17'd22884: data = 8'h16;
      17'd22885: data = 8'h1a;
      17'd22886: data = 8'h1c;
      17'd22887: data = 8'h1a;
      17'd22888: data = 8'h1b;
      17'd22889: data = 8'h1a;
      17'd22890: data = 8'h1b;
      17'd22891: data = 8'h1f;
      17'd22892: data = 8'h27;
      17'd22893: data = 8'h33;
      17'd22894: data = 8'h35;
      17'd22895: data = 8'h3d;
      17'd22896: data = 8'h45;
      17'd22897: data = 8'h47;
      17'd22898: data = 8'h4a;
      17'd22899: data = 8'h4d;
      17'd22900: data = 8'h4d;
      17'd22901: data = 8'h45;
      17'd22902: data = 8'h3c;
      17'd22903: data = 8'h2f;
      17'd22904: data = 8'h29;
      17'd22905: data = 8'h1b;
      17'd22906: data = 8'h0e;
      17'd22907: data = 8'h0a;
      17'd22908: data = 8'h05;
      17'd22909: data = 8'hfc;
      17'd22910: data = 8'hef;
      17'd22911: data = 8'heb;
      17'd22912: data = 8'he4;
      17'd22913: data = 8'he2;
      17'd22914: data = 8'he2;
      17'd22915: data = 8'he5;
      17'd22916: data = 8'he9;
      17'd22917: data = 8'he7;
      17'd22918: data = 8'hec;
      17'd22919: data = 8'hed;
      17'd22920: data = 8'heb;
      17'd22921: data = 8'hec;
      17'd22922: data = 8'hec;
      17'd22923: data = 8'hef;
      17'd22924: data = 8'hec;
      17'd22925: data = 8'he7;
      17'd22926: data = 8'he9;
      17'd22927: data = 8'he4;
      17'd22928: data = 8'he4;
      17'd22929: data = 8'he5;
      17'd22930: data = 8'heb;
      17'd22931: data = 8'hf2;
      17'd22932: data = 8'hf4;
      17'd22933: data = 8'hf4;
      17'd22934: data = 8'hfa;
      17'd22935: data = 8'hfe;
      17'd22936: data = 8'h04;
      17'd22937: data = 8'h0e;
      17'd22938: data = 8'h1c;
      17'd22939: data = 8'h27;
      17'd22940: data = 8'h2b;
      17'd22941: data = 8'h2c;
      17'd22942: data = 8'h2c;
      17'd22943: data = 8'h24;
      17'd22944: data = 8'h1e;
      17'd22945: data = 8'h1f;
      17'd22946: data = 8'h1f;
      17'd22947: data = 8'h16;
      17'd22948: data = 8'h0c;
      17'd22949: data = 8'h06;
      17'd22950: data = 8'h00;
      17'd22951: data = 8'hf9;
      17'd22952: data = 8'hf6;
      17'd22953: data = 8'hfa;
      17'd22954: data = 8'hf6;
      17'd22955: data = 8'hf6;
      17'd22956: data = 8'hf6;
      17'd22957: data = 8'hf4;
      17'd22958: data = 8'hec;
      17'd22959: data = 8'hec;
      17'd22960: data = 8'hed;
      17'd22961: data = 8'hf1;
      17'd22962: data = 8'hef;
      17'd22963: data = 8'he9;
      17'd22964: data = 8'he4;
      17'd22965: data = 8'hdb;
      17'd22966: data = 8'hd6;
      17'd22967: data = 8'hd2;
      17'd22968: data = 8'hd2;
      17'd22969: data = 8'hce;
      17'd22970: data = 8'hcb;
      17'd22971: data = 8'hca;
      17'd22972: data = 8'hc9;
      17'd22973: data = 8'hc9;
      17'd22974: data = 8'hc9;
      17'd22975: data = 8'hce;
      17'd22976: data = 8'hd6;
      17'd22977: data = 8'hdb;
      17'd22978: data = 8'he0;
      17'd22979: data = 8'he7;
      17'd22980: data = 8'he9;
      17'd22981: data = 8'heb;
      17'd22982: data = 8'hf5;
      17'd22983: data = 8'hfe;
      17'd22984: data = 8'h04;
      17'd22985: data = 8'h04;
      17'd22986: data = 8'h06;
      17'd22987: data = 8'h05;
      17'd22988: data = 8'h00;
      17'd22989: data = 8'hfe;
      17'd22990: data = 8'hfe;
      17'd22991: data = 8'h01;
      17'd22992: data = 8'h01;
      17'd22993: data = 8'hfe;
      17'd22994: data = 8'hfe;
      17'd22995: data = 8'h00;
      17'd22996: data = 8'h02;
      17'd22997: data = 8'h05;
      17'd22998: data = 8'h0d;
      17'd22999: data = 8'h12;
      17'd23000: data = 8'h15;
      17'd23001: data = 8'h19;
      17'd23002: data = 8'h13;
      17'd23003: data = 8'h13;
      17'd23004: data = 8'h11;
      17'd23005: data = 8'h11;
      17'd23006: data = 8'h0e;
      17'd23007: data = 8'h0e;
      17'd23008: data = 8'h0c;
      17'd23009: data = 8'h05;
      17'd23010: data = 8'h02;
      17'd23011: data = 8'hfe;
      17'd23012: data = 8'hfe;
      17'd23013: data = 8'hfd;
      17'd23014: data = 8'hfd;
      17'd23015: data = 8'h01;
      17'd23016: data = 8'hfd;
      17'd23017: data = 8'hf9;
      17'd23018: data = 8'hfc;
      17'd23019: data = 8'hfe;
      17'd23020: data = 8'hfc;
      17'd23021: data = 8'h05;
      17'd23022: data = 8'h09;
      17'd23023: data = 8'h06;
      17'd23024: data = 8'h0c;
      17'd23025: data = 8'h06;
      17'd23026: data = 8'h0c;
      17'd23027: data = 8'h06;
      17'd23028: data = 8'h02;
      17'd23029: data = 8'h00;
      17'd23030: data = 8'h01;
      17'd23031: data = 8'hfe;
      17'd23032: data = 8'hf5;
      17'd23033: data = 8'hfa;
      17'd23034: data = 8'hfe;
      17'd23035: data = 8'hfc;
      17'd23036: data = 8'h00;
      17'd23037: data = 8'h09;
      17'd23038: data = 8'h06;
      17'd23039: data = 8'h0c;
      17'd23040: data = 8'h15;
      17'd23041: data = 8'h1a;
      17'd23042: data = 8'h1f;
      17'd23043: data = 8'h1a;
      17'd23044: data = 8'h15;
      17'd23045: data = 8'h11;
      17'd23046: data = 8'h04;
      17'd23047: data = 8'hfa;
      17'd23048: data = 8'hf6;
      17'd23049: data = 8'hfd;
      17'd23050: data = 8'hf4;
      17'd23051: data = 8'hec;
      17'd23052: data = 8'hf6;
      17'd23053: data = 8'hec;
      17'd23054: data = 8'hec;
      17'd23055: data = 8'hf9;
      17'd23056: data = 8'h05;
      17'd23057: data = 8'h12;
      17'd23058: data = 8'h16;
      17'd23059: data = 8'h1f;
      17'd23060: data = 8'h27;
      17'd23061: data = 8'h2c;
      17'd23062: data = 8'h2f;
      17'd23063: data = 8'h43;
      17'd23064: data = 8'h45;
      17'd23065: data = 8'h3c;
      17'd23066: data = 8'h34;
      17'd23067: data = 8'h2c;
      17'd23068: data = 8'h1e;
      17'd23069: data = 8'h05;
      17'd23070: data = 8'h11;
      17'd23071: data = 8'h11;
      17'd23072: data = 8'h04;
      17'd23073: data = 8'hfc;
      17'd23074: data = 8'hf2;
      17'd23075: data = 8'hef;
      17'd23076: data = 8'he3;
      17'd23077: data = 8'he7;
      17'd23078: data = 8'hef;
      17'd23079: data = 8'hf5;
      17'd23080: data = 8'hf4;
      17'd23081: data = 8'hef;
      17'd23082: data = 8'hf2;
      17'd23083: data = 8'hed;
      17'd23084: data = 8'hec;
      17'd23085: data = 8'hf4;
      17'd23086: data = 8'hfa;
      17'd23087: data = 8'hef;
      17'd23088: data = 8'he3;
      17'd23089: data = 8'hd8;
      17'd23090: data = 8'hcb;
      17'd23091: data = 8'hc2;
      17'd23092: data = 8'hc0;
      17'd23093: data = 8'hc6;
      17'd23094: data = 8'hc6;
      17'd23095: data = 8'hbb;
      17'd23096: data = 8'hbb;
      17'd23097: data = 8'hb8;
      17'd23098: data = 8'hbb;
      17'd23099: data = 8'hc2;
      17'd23100: data = 8'hd1;
      17'd23101: data = 8'he7;
      17'd23102: data = 8'hed;
      17'd23103: data = 8'hf5;
      17'd23104: data = 8'h02;
      17'd23105: data = 8'h0a;
      17'd23106: data = 8'h15;
      17'd23107: data = 8'h23;
      17'd23108: data = 8'h31;
      17'd23109: data = 8'h33;
      17'd23110: data = 8'h2d;
      17'd23111: data = 8'h2c;
      17'd23112: data = 8'h2b;
      17'd23113: data = 8'h27;
      17'd23114: data = 8'h2c;
      17'd23115: data = 8'h33;
      17'd23116: data = 8'h33;
      17'd23117: data = 8'h31;
      17'd23118: data = 8'h27;
      17'd23119: data = 8'h26;
      17'd23120: data = 8'h27;
      17'd23121: data = 8'h27;
      17'd23122: data = 8'h2d;
      17'd23123: data = 8'h31;
      17'd23124: data = 8'h31;
      17'd23125: data = 8'h2f;
      17'd23126: data = 8'h27;
      17'd23127: data = 8'h19;
      17'd23128: data = 8'h22;
      17'd23129: data = 8'h2f;
      17'd23130: data = 8'h22;
      17'd23131: data = 8'h13;
      17'd23132: data = 8'h0d;
      17'd23133: data = 8'h01;
      17'd23134: data = 8'hf6;
      17'd23135: data = 8'hf2;
      17'd23136: data = 8'hf6;
      17'd23137: data = 8'hf2;
      17'd23138: data = 8'he7;
      17'd23139: data = 8'hdc;
      17'd23140: data = 8'hd1;
      17'd23141: data = 8'hd2;
      17'd23142: data = 8'hd8;
      17'd23143: data = 8'hd6;
      17'd23144: data = 8'hd8;
      17'd23145: data = 8'hde;
      17'd23146: data = 8'hdc;
      17'd23147: data = 8'he0;
      17'd23148: data = 8'he5;
      17'd23149: data = 8'hef;
      17'd23150: data = 8'hfd;
      17'd23151: data = 8'hfd;
      17'd23152: data = 8'hfe;
      17'd23153: data = 8'h0a;
      17'd23154: data = 8'h0d;
      17'd23155: data = 8'h0c;
      17'd23156: data = 8'h09;
      17'd23157: data = 8'h0e;
      17'd23158: data = 8'h15;
      17'd23159: data = 8'h0e;
      17'd23160: data = 8'h0d;
      17'd23161: data = 8'h0e;
      17'd23162: data = 8'h0d;
      17'd23163: data = 8'h09;
      17'd23164: data = 8'h0c;
      17'd23165: data = 8'h0d;
      17'd23166: data = 8'h11;
      17'd23167: data = 8'h13;
      17'd23168: data = 8'h13;
      17'd23169: data = 8'h13;
      17'd23170: data = 8'h1a;
      17'd23171: data = 8'h19;
      17'd23172: data = 8'h15;
      17'd23173: data = 8'h1b;
      17'd23174: data = 8'h19;
      17'd23175: data = 8'h0d;
      17'd23176: data = 8'h04;
      17'd23177: data = 8'hfe;
      17'd23178: data = 8'hfd;
      17'd23179: data = 8'hf5;
      17'd23180: data = 8'hed;
      17'd23181: data = 8'he7;
      17'd23182: data = 8'hda;
      17'd23183: data = 8'hd3;
      17'd23184: data = 8'hd3;
      17'd23185: data = 8'hd1;
      17'd23186: data = 8'hd2;
      17'd23187: data = 8'hd2;
      17'd23188: data = 8'hce;
      17'd23189: data = 8'hcd;
      17'd23190: data = 8'hd1;
      17'd23191: data = 8'hd6;
      17'd23192: data = 8'hdc;
      17'd23193: data = 8'hd8;
      17'd23194: data = 8'hda;
      17'd23195: data = 8'hde;
      17'd23196: data = 8'he0;
      17'd23197: data = 8'he3;
      17'd23198: data = 8'he4;
      17'd23199: data = 8'he9;
      17'd23200: data = 8'he2;
      17'd23201: data = 8'heb;
      17'd23202: data = 8'hdb;
      17'd23203: data = 8'he3;
      17'd23204: data = 8'hfa;
      17'd23205: data = 8'hd8;
      17'd23206: data = 8'hf4;
      17'd23207: data = 8'hfe;
      17'd23208: data = 8'hfa;
      17'd23209: data = 8'hfe;
      17'd23210: data = 8'hfe;
      17'd23211: data = 8'h16;
      17'd23212: data = 8'hfa;
      17'd23213: data = 8'h02;
      17'd23214: data = 8'h1a;
      17'd23215: data = 8'hfe;
      17'd23216: data = 8'h06;
      17'd23217: data = 8'h0d;
      17'd23218: data = 8'h0d;
      17'd23219: data = 8'h02;
      17'd23220: data = 8'h04;
      17'd23221: data = 8'h0c;
      17'd23222: data = 8'h06;
      17'd23223: data = 8'hfd;
      17'd23224: data = 8'h02;
      17'd23225: data = 8'h06;
      17'd23226: data = 8'hf9;
      17'd23227: data = 8'h0a;
      17'd23228: data = 8'h02;
      17'd23229: data = 8'hfd;
      17'd23230: data = 8'h16;
      17'd23231: data = 8'h05;
      17'd23232: data = 8'hfd;
      17'd23233: data = 8'h0a;
      17'd23234: data = 8'h06;
      17'd23235: data = 8'h04;
      17'd23236: data = 8'hfe;
      17'd23237: data = 8'h06;
      17'd23238: data = 8'h04;
      17'd23239: data = 8'hfa;
      17'd23240: data = 8'h00;
      17'd23241: data = 8'hfc;
      17'd23242: data = 8'hf6;
      17'd23243: data = 8'h06;
      17'd23244: data = 8'h04;
      17'd23245: data = 8'hf2;
      17'd23246: data = 8'h00;
      17'd23247: data = 8'h0a;
      17'd23248: data = 8'h01;
      17'd23249: data = 8'hfa;
      17'd23250: data = 8'h05;
      17'd23251: data = 8'h0e;
      17'd23252: data = 8'hfe;
      17'd23253: data = 8'h01;
      17'd23254: data = 8'h06;
      17'd23255: data = 8'h05;
      17'd23256: data = 8'h02;
      17'd23257: data = 8'h06;
      17'd23258: data = 8'h0d;
      17'd23259: data = 8'h0c;
      17'd23260: data = 8'h0d;
      17'd23261: data = 8'h02;
      17'd23262: data = 8'h04;
      17'd23263: data = 8'h0a;
      17'd23264: data = 8'h06;
      17'd23265: data = 8'h09;
      17'd23266: data = 8'h12;
      17'd23267: data = 8'h1b;
      17'd23268: data = 8'h1a;
      17'd23269: data = 8'h1a;
      17'd23270: data = 8'h13;
      17'd23271: data = 8'h05;
      17'd23272: data = 8'h01;
      17'd23273: data = 8'hfa;
      17'd23274: data = 8'hf1;
      17'd23275: data = 8'he9;
      17'd23276: data = 8'hef;
      17'd23277: data = 8'heb;
      17'd23278: data = 8'he2;
      17'd23279: data = 8'hed;
      17'd23280: data = 8'hf2;
      17'd23281: data = 8'hf2;
      17'd23282: data = 8'hfd;
      17'd23283: data = 8'h09;
      17'd23284: data = 8'h0e;
      17'd23285: data = 8'h12;
      17'd23286: data = 8'h1a;
      17'd23287: data = 8'h24;
      17'd23288: data = 8'h2f;
      17'd23289: data = 8'h35;
      17'd23290: data = 8'h3d;
      17'd23291: data = 8'h3a;
      17'd23292: data = 8'h33;
      17'd23293: data = 8'h29;
      17'd23294: data = 8'h1e;
      17'd23295: data = 8'h1e;
      17'd23296: data = 8'h19;
      17'd23297: data = 8'h13;
      17'd23298: data = 8'h0d;
      17'd23299: data = 8'h01;
      17'd23300: data = 8'hfa;
      17'd23301: data = 8'hf1;
      17'd23302: data = 8'hef;
      17'd23303: data = 8'hf2;
      17'd23304: data = 8'hef;
      17'd23305: data = 8'hed;
      17'd23306: data = 8'hed;
      17'd23307: data = 8'hef;
      17'd23308: data = 8'hed;
      17'd23309: data = 8'hed;
      17'd23310: data = 8'hf2;
      17'd23311: data = 8'hf2;
      17'd23312: data = 8'hed;
      17'd23313: data = 8'hec;
      17'd23314: data = 8'he3;
      17'd23315: data = 8'hd8;
      17'd23316: data = 8'hd3;
      17'd23317: data = 8'hd3;
      17'd23318: data = 8'hd1;
      17'd23319: data = 8'hce;
      17'd23320: data = 8'hcb;
      17'd23321: data = 8'hcb;
      17'd23322: data = 8'hca;
      17'd23323: data = 8'hc6;
      17'd23324: data = 8'hcb;
      17'd23325: data = 8'hcd;
      17'd23326: data = 8'hce;
      17'd23327: data = 8'hd5;
      17'd23328: data = 8'he2;
      17'd23329: data = 8'hed;
      17'd23330: data = 8'hf4;
      17'd23331: data = 8'hfe;
      17'd23332: data = 8'h0a;
      17'd23333: data = 8'h11;
      17'd23334: data = 8'h1a;
      17'd23335: data = 8'h23;
      17'd23336: data = 8'h2b;
      17'd23337: data = 8'h31;
      17'd23338: data = 8'h35;
      17'd23339: data = 8'h39;
      17'd23340: data = 8'h3a;
      17'd23341: data = 8'h3c;
      17'd23342: data = 8'h3a;
      17'd23343: data = 8'h3c;
      17'd23344: data = 8'h36;
      17'd23345: data = 8'h31;
      17'd23346: data = 8'h27;
      17'd23347: data = 8'h22;
      17'd23348: data = 8'h1c;
      17'd23349: data = 8'h1a;
      17'd23350: data = 8'h1b;
      17'd23351: data = 8'h1b;
      17'd23352: data = 8'h1a;
      17'd23353: data = 8'h16;
      17'd23354: data = 8'h13;
      17'd23355: data = 8'h11;
      17'd23356: data = 8'h11;
      17'd23357: data = 8'h11;
      17'd23358: data = 8'h0e;
      17'd23359: data = 8'h0d;
      17'd23360: data = 8'h09;
      17'd23361: data = 8'h05;
      17'd23362: data = 8'h02;
      17'd23363: data = 8'h00;
      17'd23364: data = 8'hfa;
      17'd23365: data = 8'hf4;
      17'd23366: data = 8'hef;
      17'd23367: data = 8'he4;
      17'd23368: data = 8'hdc;
      17'd23369: data = 8'hdc;
      17'd23370: data = 8'hda;
      17'd23371: data = 8'hd8;
      17'd23372: data = 8'hda;
      17'd23373: data = 8'hde;
      17'd23374: data = 8'he2;
      17'd23375: data = 8'he4;
      17'd23376: data = 8'hed;
      17'd23377: data = 8'hf2;
      17'd23378: data = 8'hfa;
      17'd23379: data = 8'h04;
      17'd23380: data = 8'h0a;
      17'd23381: data = 8'h11;
      17'd23382: data = 8'h15;
      17'd23383: data = 8'h1b;
      17'd23384: data = 8'h1c;
      17'd23385: data = 8'h1a;
      17'd23386: data = 8'h16;
      17'd23387: data = 8'h16;
      17'd23388: data = 8'h15;
      17'd23389: data = 8'h11;
      17'd23390: data = 8'h12;
      17'd23391: data = 8'h11;
      17'd23392: data = 8'h0e;
      17'd23393: data = 8'h0c;
      17'd23394: data = 8'h0c;
      17'd23395: data = 8'h0c;
      17'd23396: data = 8'h09;
      17'd23397: data = 8'h06;
      17'd23398: data = 8'h05;
      17'd23399: data = 8'h06;
      17'd23400: data = 8'h05;
      17'd23401: data = 8'h02;
      17'd23402: data = 8'h01;
      17'd23403: data = 8'hfd;
      17'd23404: data = 8'hfc;
      17'd23405: data = 8'hfa;
      17'd23406: data = 8'hf5;
      17'd23407: data = 8'hf1;
      17'd23408: data = 8'heb;
      17'd23409: data = 8'he7;
      17'd23410: data = 8'he3;
      17'd23411: data = 8'hde;
      17'd23412: data = 8'hdc;
      17'd23413: data = 8'hdb;
      17'd23414: data = 8'hd8;
      17'd23415: data = 8'hd5;
      17'd23416: data = 8'hd5;
      17'd23417: data = 8'hd3;
      17'd23418: data = 8'hd5;
      17'd23419: data = 8'hd6;
      17'd23420: data = 8'hd8;
      17'd23421: data = 8'hda;
      17'd23422: data = 8'hdc;
      17'd23423: data = 8'he2;
      17'd23424: data = 8'he4;
      17'd23425: data = 8'heb;
      17'd23426: data = 8'hed;
      17'd23427: data = 8'hf1;
      17'd23428: data = 8'hf5;
      17'd23429: data = 8'hf6;
      17'd23430: data = 8'hf6;
      17'd23431: data = 8'hfd;
      17'd23432: data = 8'h00;
      17'd23433: data = 8'h00;
      17'd23434: data = 8'h01;
      17'd23435: data = 8'h02;
      17'd23436: data = 8'h00;
      17'd23437: data = 8'hfe;
      17'd23438: data = 8'h00;
      17'd23439: data = 8'h00;
      17'd23440: data = 8'hfd;
      17'd23441: data = 8'hfc;
      17'd23442: data = 8'hfc;
      17'd23443: data = 8'hf6;
      17'd23444: data = 8'hf5;
      17'd23445: data = 8'hf6;
      17'd23446: data = 8'hf9;
      17'd23447: data = 8'hfc;
      17'd23448: data = 8'h00;
      17'd23449: data = 8'h02;
      17'd23450: data = 8'h05;
      17'd23451: data = 8'h0a;
      17'd23452: data = 8'h0c;
      17'd23453: data = 8'h0d;
      17'd23454: data = 8'h0d;
      17'd23455: data = 8'h0e;
      17'd23456: data = 8'h0c;
      17'd23457: data = 8'h04;
      17'd23458: data = 8'h04;
      17'd23459: data = 8'h00;
      17'd23460: data = 8'hfd;
      17'd23461: data = 8'hfa;
      17'd23462: data = 8'hfc;
      17'd23463: data = 8'hfa;
      17'd23464: data = 8'hfc;
      17'd23465: data = 8'hfe;
      17'd23466: data = 8'h00;
      17'd23467: data = 8'h02;
      17'd23468: data = 8'h04;
      17'd23469: data = 8'h05;
      17'd23470: data = 8'h05;
      17'd23471: data = 8'h06;
      17'd23472: data = 8'h09;
      17'd23473: data = 8'h06;
      17'd23474: data = 8'h0a;
      17'd23475: data = 8'h0c;
      17'd23476: data = 8'h0c;
      17'd23477: data = 8'h09;
      17'd23478: data = 8'h04;
      17'd23479: data = 8'h04;
      17'd23480: data = 8'h05;
      17'd23481: data = 8'h02;
      17'd23482: data = 8'h01;
      17'd23483: data = 8'h00;
      17'd23484: data = 8'h00;
      17'd23485: data = 8'h04;
      17'd23486: data = 8'h02;
      17'd23487: data = 8'h05;
      17'd23488: data = 8'h04;
      17'd23489: data = 8'h09;
      17'd23490: data = 8'h06;
      17'd23491: data = 8'h05;
      17'd23492: data = 8'h0a;
      17'd23493: data = 8'h0a;
      17'd23494: data = 8'h0e;
      17'd23495: data = 8'h0d;
      17'd23496: data = 8'h16;
      17'd23497: data = 8'h15;
      17'd23498: data = 8'h0e;
      17'd23499: data = 8'h0a;
      17'd23500: data = 8'h00;
      17'd23501: data = 8'hfd;
      17'd23502: data = 8'hf4;
      17'd23503: data = 8'hf1;
      17'd23504: data = 8'hef;
      17'd23505: data = 8'hef;
      17'd23506: data = 8'hed;
      17'd23507: data = 8'he9;
      17'd23508: data = 8'hec;
      17'd23509: data = 8'he9;
      17'd23510: data = 8'hf2;
      17'd23511: data = 8'hfd;
      17'd23512: data = 8'h05;
      17'd23513: data = 8'h0c;
      17'd23514: data = 8'h11;
      17'd23515: data = 8'h1b;
      17'd23516: data = 8'h22;
      17'd23517: data = 8'h2b;
      17'd23518: data = 8'h33;
      17'd23519: data = 8'h39;
      17'd23520: data = 8'h35;
      17'd23521: data = 8'h2f;
      17'd23522: data = 8'h2c;
      17'd23523: data = 8'h27;
      17'd23524: data = 8'h26;
      17'd23525: data = 8'h1f;
      17'd23526: data = 8'h1e;
      17'd23527: data = 8'h15;
      17'd23528: data = 8'h09;
      17'd23529: data = 8'h02;
      17'd23530: data = 8'hfa;
      17'd23531: data = 8'hf4;
      17'd23532: data = 8'hed;
      17'd23533: data = 8'he9;
      17'd23534: data = 8'he4;
      17'd23535: data = 8'he3;
      17'd23536: data = 8'hdc;
      17'd23537: data = 8'hdc;
      17'd23538: data = 8'he0;
      17'd23539: data = 8'he4;
      17'd23540: data = 8'he5;
      17'd23541: data = 8'heb;
      17'd23542: data = 8'hed;
      17'd23543: data = 8'he9;
      17'd23544: data = 8'he9;
      17'd23545: data = 8'heb;
      17'd23546: data = 8'heb;
      17'd23547: data = 8'he7;
      17'd23548: data = 8'he3;
      17'd23549: data = 8'he4;
      17'd23550: data = 8'hde;
      17'd23551: data = 8'hd3;
      17'd23552: data = 8'hce;
      17'd23553: data = 8'hce;
      17'd23554: data = 8'hce;
      17'd23555: data = 8'hce;
      17'd23556: data = 8'hd8;
      17'd23557: data = 8'hdb;
      17'd23558: data = 8'he2;
      17'd23559: data = 8'he9;
      17'd23560: data = 8'hf4;
      17'd23561: data = 8'h01;
      17'd23562: data = 8'h0c;
      17'd23563: data = 8'h1a;
      17'd23564: data = 8'h26;
      17'd23565: data = 8'h2d;
      17'd23566: data = 8'h33;
      17'd23567: data = 8'h3a;
      17'd23568: data = 8'h3d;
      17'd23569: data = 8'h3d;
      17'd23570: data = 8'h3e;
      17'd23571: data = 8'h3d;
      17'd23572: data = 8'h3a;
      17'd23573: data = 8'h33;
      17'd23574: data = 8'h2b;
      17'd23575: data = 8'h27;
      17'd23576: data = 8'h23;
      17'd23577: data = 8'h1b;
      17'd23578: data = 8'h16;
      17'd23579: data = 8'h12;
      17'd23580: data = 8'h0e;
      17'd23581: data = 8'h0a;
      17'd23582: data = 8'h04;
      17'd23583: data = 8'h02;
      17'd23584: data = 8'h02;
      17'd23585: data = 8'h04;
      17'd23586: data = 8'h02;
      17'd23587: data = 8'h02;
      17'd23588: data = 8'h01;
      17'd23589: data = 8'h00;
      17'd23590: data = 8'h01;
      17'd23591: data = 8'h00;
      17'd23592: data = 8'hfd;
      17'd23593: data = 8'hfd;
      17'd23594: data = 8'hfd;
      17'd23595: data = 8'hf9;
      17'd23596: data = 8'hf4;
      17'd23597: data = 8'hed;
      17'd23598: data = 8'heb;
      17'd23599: data = 8'he9;
      17'd23600: data = 8'he5;
      17'd23601: data = 8'he4;
      17'd23602: data = 8'he3;
      17'd23603: data = 8'he2;
      17'd23604: data = 8'he2;
      17'd23605: data = 8'he4;
      17'd23606: data = 8'he7;
      17'd23607: data = 8'hec;
      17'd23608: data = 8'hf2;
      17'd23609: data = 8'hf9;
      17'd23610: data = 8'hfe;
      17'd23611: data = 8'h05;
      17'd23612: data = 8'h0e;
      17'd23613: data = 8'h19;
      17'd23614: data = 8'h19;
      17'd23615: data = 8'h11;
      17'd23616: data = 8'h19;
      17'd23617: data = 8'h22;
      17'd23618: data = 8'h1c;
      17'd23619: data = 8'h1e;
      17'd23620: data = 8'h24;
      17'd23621: data = 8'h22;
      17'd23622: data = 8'h15;
      17'd23623: data = 8'h11;
      17'd23624: data = 8'h0c;
      17'd23625: data = 8'h02;
      17'd23626: data = 8'hfe;
      17'd23627: data = 8'hfe;
      17'd23628: data = 8'hf6;
      17'd23629: data = 8'hed;
      17'd23630: data = 8'hef;
      17'd23631: data = 8'hf2;
      17'd23632: data = 8'hed;
      17'd23633: data = 8'heb;
      17'd23634: data = 8'hf2;
      17'd23635: data = 8'hf1;
      17'd23636: data = 8'he9;
      17'd23637: data = 8'hf1;
      17'd23638: data = 8'hfc;
      17'd23639: data = 8'hf9;
      17'd23640: data = 8'hf5;
      17'd23641: data = 8'hf5;
      17'd23642: data = 8'hef;
      17'd23643: data = 8'hec;
      17'd23644: data = 8'he9;
      17'd23645: data = 8'he0;
      17'd23646: data = 8'hdb;
      17'd23647: data = 8'hde;
      17'd23648: data = 8'hda;
      17'd23649: data = 8'hd8;
      17'd23650: data = 8'hdc;
      17'd23651: data = 8'hdb;
      17'd23652: data = 8'hda;
      17'd23653: data = 8'hde;
      17'd23654: data = 8'he7;
      17'd23655: data = 8'he7;
      17'd23656: data = 8'he4;
      17'd23657: data = 8'hed;
      17'd23658: data = 8'hf9;
      17'd23659: data = 8'hf5;
      17'd23660: data = 8'hf5;
      17'd23661: data = 8'hfe;
      17'd23662: data = 8'h02;
      17'd23663: data = 8'hfa;
      17'd23664: data = 8'hfc;
      17'd23665: data = 8'h02;
      17'd23666: data = 8'hfc;
      17'd23667: data = 8'hf5;
      17'd23668: data = 8'hfd;
      17'd23669: data = 8'h01;
      17'd23670: data = 8'hfa;
      17'd23671: data = 8'hf9;
      17'd23672: data = 8'hfa;
      17'd23673: data = 8'hf9;
      17'd23674: data = 8'hf4;
      17'd23675: data = 8'hf6;
      17'd23676: data = 8'hfc;
      17'd23677: data = 8'hfc;
      17'd23678: data = 8'hfd;
      17'd23679: data = 8'h00;
      17'd23680: data = 8'h02;
      17'd23681: data = 8'h02;
      17'd23682: data = 8'h05;
      17'd23683: data = 8'h0c;
      17'd23684: data = 8'h0c;
      17'd23685: data = 8'h09;
      17'd23686: data = 8'h0c;
      17'd23687: data = 8'h0e;
      17'd23688: data = 8'h0d;
      17'd23689: data = 8'h0a;
      17'd23690: data = 8'h0d;
      17'd23691: data = 8'h0c;
      17'd23692: data = 8'h06;
      17'd23693: data = 8'h05;
      17'd23694: data = 8'h02;
      17'd23695: data = 8'h00;
      17'd23696: data = 8'hfd;
      17'd23697: data = 8'hfd;
      17'd23698: data = 8'hfe;
      17'd23699: data = 8'hfc;
      17'd23700: data = 8'hf6;
      17'd23701: data = 8'hf9;
      17'd23702: data = 8'hfe;
      17'd23703: data = 8'hfc;
      17'd23704: data = 8'hfd;
      17'd23705: data = 8'h01;
      17'd23706: data = 8'h04;
      17'd23707: data = 8'h04;
      17'd23708: data = 8'h06;
      17'd23709: data = 8'h0a;
      17'd23710: data = 8'h0a;
      17'd23711: data = 8'h0a;
      17'd23712: data = 8'h0d;
      17'd23713: data = 8'h0c;
      17'd23714: data = 8'h09;
      17'd23715: data = 8'h02;
      17'd23716: data = 8'h02;
      17'd23717: data = 8'h01;
      17'd23718: data = 8'hfd;
      17'd23719: data = 8'hfc;
      17'd23720: data = 8'hfe;
      17'd23721: data = 8'hfe;
      17'd23722: data = 8'hfd;
      17'd23723: data = 8'h02;
      17'd23724: data = 8'h09;
      17'd23725: data = 8'h09;
      17'd23726: data = 8'h0d;
      17'd23727: data = 8'h12;
      17'd23728: data = 8'h0e;
      17'd23729: data = 8'h05;
      17'd23730: data = 8'h02;
      17'd23731: data = 8'h04;
      17'd23732: data = 8'h02;
      17'd23733: data = 8'h00;
      17'd23734: data = 8'h01;
      17'd23735: data = 8'hfe;
      17'd23736: data = 8'hf5;
      17'd23737: data = 8'hf2;
      17'd23738: data = 8'hf4;
      17'd23739: data = 8'hf1;
      17'd23740: data = 8'hf5;
      17'd23741: data = 8'hfd;
      17'd23742: data = 8'hfe;
      17'd23743: data = 8'h00;
      17'd23744: data = 8'h0a;
      17'd23745: data = 8'h15;
      17'd23746: data = 8'h15;
      17'd23747: data = 8'h22;
      17'd23748: data = 8'h2c;
      17'd23749: data = 8'h2b;
      17'd23750: data = 8'h27;
      17'd23751: data = 8'h2f;
      17'd23752: data = 8'h31;
      17'd23753: data = 8'h27;
      17'd23754: data = 8'h27;
      17'd23755: data = 8'h26;
      17'd23756: data = 8'h1c;
      17'd23757: data = 8'h0e;
      17'd23758: data = 8'h09;
      17'd23759: data = 8'h01;
      17'd23760: data = 8'hf6;
      17'd23761: data = 8'hf4;
      17'd23762: data = 8'hf1;
      17'd23763: data = 8'hec;
      17'd23764: data = 8'heb;
      17'd23765: data = 8'he5;
      17'd23766: data = 8'hde;
      17'd23767: data = 8'hdb;
      17'd23768: data = 8'he0;
      17'd23769: data = 8'hde;
      17'd23770: data = 8'hda;
      17'd23771: data = 8'hde;
      17'd23772: data = 8'he4;
      17'd23773: data = 8'he0;
      17'd23774: data = 8'hde;
      17'd23775: data = 8'he7;
      17'd23776: data = 8'he9;
      17'd23777: data = 8'he4;
      17'd23778: data = 8'he7;
      17'd23779: data = 8'heb;
      17'd23780: data = 8'he4;
      17'd23781: data = 8'hde;
      17'd23782: data = 8'he4;
      17'd23783: data = 8'he9;
      17'd23784: data = 8'he4;
      17'd23785: data = 8'he7;
      17'd23786: data = 8'hed;
      17'd23787: data = 8'hed;
      17'd23788: data = 8'heb;
      17'd23789: data = 8'hed;
      17'd23790: data = 8'hf5;
      17'd23791: data = 8'hfa;
      17'd23792: data = 8'hfd;
      17'd23793: data = 8'h05;
      17'd23794: data = 8'h0e;
      17'd23795: data = 8'h13;
      17'd23796: data = 8'h19;
      17'd23797: data = 8'h24;
      17'd23798: data = 8'h2c;
      17'd23799: data = 8'h2f;
      17'd23800: data = 8'h35;
      17'd23801: data = 8'h3a;
      17'd23802: data = 8'h3c;
      17'd23803: data = 8'h3c;
      17'd23804: data = 8'h3c;
      17'd23805: data = 8'h39;
      17'd23806: data = 8'h31;
      17'd23807: data = 8'h2c;
      17'd23808: data = 8'h26;
      17'd23809: data = 8'h1e;
      17'd23810: data = 8'h15;
      17'd23811: data = 8'h0c;
      17'd23812: data = 8'h06;
      17'd23813: data = 8'h02;
      17'd23814: data = 8'hfe;
      17'd23815: data = 8'hfa;
      17'd23816: data = 8'hf6;
      17'd23817: data = 8'hf5;
      17'd23818: data = 8'hf2;
      17'd23819: data = 8'hf1;
      17'd23820: data = 8'hf2;
      17'd23821: data = 8'hf4;
      17'd23822: data = 8'hf5;
      17'd23823: data = 8'hf6;
      17'd23824: data = 8'hf9;
      17'd23825: data = 8'hf5;
      17'd23826: data = 8'hf5;
      17'd23827: data = 8'hf4;
      17'd23828: data = 8'hf4;
      17'd23829: data = 8'hf4;
      17'd23830: data = 8'hf4;
      17'd23831: data = 8'hf1;
      17'd23832: data = 8'hef;
      17'd23833: data = 8'hf1;
      17'd23834: data = 8'hef;
      17'd23835: data = 8'hf2;
      17'd23836: data = 8'hf2;
      17'd23837: data = 8'hf2;
      17'd23838: data = 8'hf4;
      17'd23839: data = 8'hf5;
      17'd23840: data = 8'hfa;
      17'd23841: data = 8'hfc;
      17'd23842: data = 8'h00;
      17'd23843: data = 8'h06;
      17'd23844: data = 8'h0a;
      17'd23845: data = 8'h11;
      17'd23846: data = 8'h11;
      17'd23847: data = 8'h05;
      17'd23848: data = 8'h0a;
      17'd23849: data = 8'h1a;
      17'd23850: data = 8'h19;
      17'd23851: data = 8'h12;
      17'd23852: data = 8'h1e;
      17'd23853: data = 8'h23;
      17'd23854: data = 8'h11;
      17'd23855: data = 8'h0a;
      17'd23856: data = 8'h0d;
      17'd23857: data = 8'h04;
      17'd23858: data = 8'hfd;
      17'd23859: data = 8'h01;
      17'd23860: data = 8'h00;
      17'd23861: data = 8'hf5;
      17'd23862: data = 8'hf5;
      17'd23863: data = 8'hfc;
      17'd23864: data = 8'hf4;
      17'd23865: data = 8'heb;
      17'd23866: data = 8'hec;
      17'd23867: data = 8'heb;
      17'd23868: data = 8'he0;
      17'd23869: data = 8'he2;
      17'd23870: data = 8'hec;
      17'd23871: data = 8'hf1;
      17'd23872: data = 8'heb;
      17'd23873: data = 8'hec;
      17'd23874: data = 8'hf1;
      17'd23875: data = 8'heb;
      17'd23876: data = 8'he4;
      17'd23877: data = 8'he3;
      17'd23878: data = 8'he3;
      17'd23879: data = 8'he4;
      17'd23880: data = 8'he3;
      17'd23881: data = 8'he3;
      17'd23882: data = 8'he5;
      17'd23883: data = 8'hde;
      17'd23884: data = 8'hda;
      17'd23885: data = 8'hdb;
      17'd23886: data = 8'he2;
      17'd23887: data = 8'he0;
      17'd23888: data = 8'hdb;
      17'd23889: data = 8'he7;
      17'd23890: data = 8'hf1;
      17'd23891: data = 8'hec;
      17'd23892: data = 8'hef;
      17'd23893: data = 8'hfc;
      17'd23894: data = 8'hfd;
      17'd23895: data = 8'hf6;
      17'd23896: data = 8'hfd;
      17'd23897: data = 8'h05;
      17'd23898: data = 8'h02;
      17'd23899: data = 8'hfd;
      17'd23900: data = 8'h05;
      17'd23901: data = 8'h09;
      17'd23902: data = 8'hfa;
      17'd23903: data = 8'hf5;
      17'd23904: data = 8'hfc;
      17'd23905: data = 8'hf9;
      17'd23906: data = 8'hf4;
      17'd23907: data = 8'hf9;
      17'd23908: data = 8'hfd;
      17'd23909: data = 8'hfd;
      17'd23910: data = 8'h00;
      17'd23911: data = 8'h09;
      17'd23912: data = 8'h0d;
      17'd23913: data = 8'h0d;
      17'd23914: data = 8'h11;
      17'd23915: data = 8'h13;
      17'd23916: data = 8'h0e;
      17'd23917: data = 8'h0d;
      17'd23918: data = 8'h12;
      17'd23919: data = 8'h0d;
      17'd23920: data = 8'h06;
      17'd23921: data = 8'h04;
      17'd23922: data = 8'h02;
      17'd23923: data = 8'h01;
      17'd23924: data = 8'hfe;
      17'd23925: data = 8'hfe;
      17'd23926: data = 8'hfe;
      17'd23927: data = 8'hfd;
      17'd23928: data = 8'h00;
      17'd23929: data = 8'h00;
      17'd23930: data = 8'hfc;
      17'd23931: data = 8'hfc;
      17'd23932: data = 8'hfe;
      17'd23933: data = 8'hfd;
      17'd23934: data = 8'hfa;
      17'd23935: data = 8'hfd;
      17'd23936: data = 8'h00;
      17'd23937: data = 8'hfd;
      17'd23938: data = 8'hfe;
      17'd23939: data = 8'h02;
      17'd23940: data = 8'h00;
      17'd23941: data = 8'h00;
      17'd23942: data = 8'h02;
      17'd23943: data = 8'h02;
      17'd23944: data = 8'h02;
      17'd23945: data = 8'h02;
      17'd23946: data = 8'h04;
      17'd23947: data = 8'h06;
      17'd23948: data = 8'h09;
      17'd23949: data = 8'h0c;
      17'd23950: data = 8'h0c;
      17'd23951: data = 8'h06;
      17'd23952: data = 8'h09;
      17'd23953: data = 8'h09;
      17'd23954: data = 8'h0a;
      17'd23955: data = 8'h0d;
      17'd23956: data = 8'h11;
      17'd23957: data = 8'h15;
      17'd23958: data = 8'h13;
      17'd23959: data = 8'h0c;
      17'd23960: data = 8'h04;
      17'd23961: data = 8'h04;
      17'd23962: data = 8'h04;
      17'd23963: data = 8'hfd;
      17'd23964: data = 8'hfd;
      17'd23965: data = 8'h00;
      17'd23966: data = 8'hfc;
      17'd23967: data = 8'hf6;
      17'd23968: data = 8'hfc;
      17'd23969: data = 8'hfe;
      17'd23970: data = 8'hfc;
      17'd23971: data = 8'h02;
      17'd23972: data = 8'h09;
      17'd23973: data = 8'h09;
      17'd23974: data = 8'h05;
      17'd23975: data = 8'h0d;
      17'd23976: data = 8'h12;
      17'd23977: data = 8'h11;
      17'd23978: data = 8'h13;
      17'd23979: data = 8'h1c;
      17'd23980: data = 8'h1e;
      17'd23981: data = 8'h1b;
      17'd23982: data = 8'h1f;
      17'd23983: data = 8'h24;
      17'd23984: data = 8'h24;
      17'd23985: data = 8'h23;
      17'd23986: data = 8'h22;
      17'd23987: data = 8'h1c;
      17'd23988: data = 8'h15;
      17'd23989: data = 8'h0c;
      17'd23990: data = 8'h01;
      17'd23991: data = 8'hfc;
      17'd23992: data = 8'hf5;
      17'd23993: data = 8'hef;
      17'd23994: data = 8'hec;
      17'd23995: data = 8'hec;
      17'd23996: data = 8'he4;
      17'd23997: data = 8'hdb;
      17'd23998: data = 8'hde;
      17'd23999: data = 8'he2;
      17'd24000: data = 8'hde;
      17'd24001: data = 8'he2;
      17'd24002: data = 8'he5;
      17'd24003: data = 8'he7;
      17'd24004: data = 8'he4;
      17'd24005: data = 8'he5;
      17'd24006: data = 8'hec;
      17'd24007: data = 8'hed;
      17'd24008: data = 8'hec;
      17'd24009: data = 8'hf2;
      17'd24010: data = 8'hf4;
      17'd24011: data = 8'hec;
      17'd24012: data = 8'he9;
      17'd24013: data = 8'heb;
      17'd24014: data = 8'hec;
      17'd24015: data = 8'heb;
      17'd24016: data = 8'hed;
      17'd24017: data = 8'hf4;
      17'd24018: data = 8'hf4;
      17'd24019: data = 8'hf1;
      17'd24020: data = 8'hf6;
      17'd24021: data = 8'hfd;
      17'd24022: data = 8'hfe;
      17'd24023: data = 8'h02;
      17'd24024: data = 8'h0c;
      17'd24025: data = 8'h12;
      17'd24026: data = 8'h11;
      17'd24027: data = 8'h16;
      17'd24028: data = 8'h1c;
      17'd24029: data = 8'h1e;
      17'd24030: data = 8'h23;
      17'd24031: data = 8'h2b;
      17'd24032: data = 8'h2d;
      17'd24033: data = 8'h2c;
      17'd24034: data = 8'h2d;
      17'd24035: data = 8'h2f;
      17'd24036: data = 8'h2d;
      17'd24037: data = 8'h29;
      17'd24038: data = 8'h27;
      17'd24039: data = 8'h23;
      17'd24040: data = 8'h1b;
      17'd24041: data = 8'h1a;
      17'd24042: data = 8'h15;
      17'd24043: data = 8'h0e;
      17'd24044: data = 8'h09;
      17'd24045: data = 8'h04;
      17'd24046: data = 8'hfe;
      17'd24047: data = 8'hf6;
      17'd24048: data = 8'hf1;
      17'd24049: data = 8'hec;
      17'd24050: data = 8'he7;
      17'd24051: data = 8'he4;
      17'd24052: data = 8'he5;
      17'd24053: data = 8'heb;
      17'd24054: data = 8'hec;
      17'd24055: data = 8'hef;
      17'd24056: data = 8'hf1;
      17'd24057: data = 8'hf4;
      17'd24058: data = 8'hf9;
      17'd24059: data = 8'hf9;
      17'd24060: data = 8'hfa;
      17'd24061: data = 8'hfd;
      17'd24062: data = 8'hfd;
      17'd24063: data = 8'hfc;
      17'd24064: data = 8'hfc;
      17'd24065: data = 8'hfc;
      17'd24066: data = 8'hf9;
      17'd24067: data = 8'hf6;
      17'd24068: data = 8'hf9;
      17'd24069: data = 8'hf9;
      17'd24070: data = 8'hfa;
      17'd24071: data = 8'hfc;
      17'd24072: data = 8'hfd;
      17'd24073: data = 8'hfe;
      17'd24074: data = 8'h01;
      17'd24075: data = 8'h04;
      17'd24076: data = 8'h05;
      17'd24077: data = 8'h09;
      17'd24078: data = 8'h0a;
      17'd24079: data = 8'h0c;
      17'd24080: data = 8'h11;
      17'd24081: data = 8'h12;
      17'd24082: data = 8'h13;
      17'd24083: data = 8'h19;
      17'd24084: data = 8'h19;
      17'd24085: data = 8'h15;
      17'd24086: data = 8'h11;
      17'd24087: data = 8'h0e;
      17'd24088: data = 8'h09;
      17'd24089: data = 8'h06;
      17'd24090: data = 8'h04;
      17'd24091: data = 8'h00;
      17'd24092: data = 8'hfc;
      17'd24093: data = 8'hf9;
      17'd24094: data = 8'hf5;
      17'd24095: data = 8'hf4;
      17'd24096: data = 8'hef;
      17'd24097: data = 8'hec;
      17'd24098: data = 8'heb;
      17'd24099: data = 8'he7;
      17'd24100: data = 8'he5;
      17'd24101: data = 8'he4;
      17'd24102: data = 8'he3;
      17'd24103: data = 8'he3;
      17'd24104: data = 8'he4;
      17'd24105: data = 8'he0;
      17'd24106: data = 8'he0;
      17'd24107: data = 8'he2;
      17'd24108: data = 8'he0;
      17'd24109: data = 8'he0;
      17'd24110: data = 8'he2;
      17'd24111: data = 8'he3;
      17'd24112: data = 8'he3;
      17'd24113: data = 8'he3;
      17'd24114: data = 8'he7;
      17'd24115: data = 8'he9;
      17'd24116: data = 8'he9;
      17'd24117: data = 8'hed;
      17'd24118: data = 8'hed;
      17'd24119: data = 8'hed;
      17'd24120: data = 8'hef;
      17'd24121: data = 8'hef;
      17'd24122: data = 8'hef;
      17'd24123: data = 8'hed;
      17'd24124: data = 8'hed;
      17'd24125: data = 8'hf1;
      17'd24126: data = 8'hf2;
      17'd24127: data = 8'hf4;
      17'd24128: data = 8'hf9;
      17'd24129: data = 8'hfa;
      17'd24130: data = 8'hfc;
      17'd24131: data = 8'hfe;
      17'd24132: data = 8'h00;
      17'd24133: data = 8'h00;
      17'd24134: data = 8'h01;
      17'd24135: data = 8'h04;
      17'd24136: data = 8'h05;
      17'd24137: data = 8'h05;
      17'd24138: data = 8'h04;
      17'd24139: data = 8'h04;
      17'd24140: data = 8'h05;
      17'd24141: data = 8'h05;
      17'd24142: data = 8'h06;
      17'd24143: data = 8'h09;
      17'd24144: data = 8'h09;
      17'd24145: data = 8'h09;
      17'd24146: data = 8'h05;
      17'd24147: data = 8'h04;
      17'd24148: data = 8'h06;
      17'd24149: data = 8'h05;
      17'd24150: data = 8'h04;
      17'd24151: data = 8'h05;
      17'd24152: data = 8'h04;
      17'd24153: data = 8'h01;
      17'd24154: data = 8'h02;
      17'd24155: data = 8'h02;
      17'd24156: data = 8'h00;
      17'd24157: data = 8'h00;
      17'd24158: data = 8'h01;
      17'd24159: data = 8'hfc;
      17'd24160: data = 8'hf6;
      17'd24161: data = 8'hf9;
      17'd24162: data = 8'hf6;
      17'd24163: data = 8'hf4;
      17'd24164: data = 8'hf5;
      17'd24165: data = 8'hfc;
      17'd24166: data = 8'hfc;
      17'd24167: data = 8'hfc;
      17'd24168: data = 8'h02;
      17'd24169: data = 8'h05;
      17'd24170: data = 8'h06;
      17'd24171: data = 8'h09;
      17'd24172: data = 8'h0d;
      17'd24173: data = 8'h12;
      17'd24174: data = 8'h11;
      17'd24175: data = 8'h11;
      17'd24176: data = 8'h12;
      17'd24177: data = 8'h11;
      17'd24178: data = 8'h0a;
      17'd24179: data = 8'h0a;
      17'd24180: data = 8'h0d;
      17'd24181: data = 8'h09;
      17'd24182: data = 8'h02;
      17'd24183: data = 8'h09;
      17'd24184: data = 8'h09;
      17'd24185: data = 8'h05;
      17'd24186: data = 8'h09;
      17'd24187: data = 8'h11;
      17'd24188: data = 8'h13;
      17'd24189: data = 8'h13;
      17'd24190: data = 8'h16;
      17'd24191: data = 8'h19;
      17'd24192: data = 8'h0d;
      17'd24193: data = 8'h01;
      17'd24194: data = 8'h04;
      17'd24195: data = 8'h01;
      17'd24196: data = 8'hfa;
      17'd24197: data = 8'hfa;
      17'd24198: data = 8'hfc;
      17'd24199: data = 8'hf4;
      17'd24200: data = 8'hef;
      17'd24201: data = 8'hf5;
      17'd24202: data = 8'hf4;
      17'd24203: data = 8'hf5;
      17'd24204: data = 8'hfd;
      17'd24205: data = 8'h02;
      17'd24206: data = 8'h05;
      17'd24207: data = 8'h05;
      17'd24208: data = 8'h0a;
      17'd24209: data = 8'h0e;
      17'd24210: data = 8'h13;
      17'd24211: data = 8'h19;
      17'd24212: data = 8'h19;
      17'd24213: data = 8'h1b;
      17'd24214: data = 8'h1c;
      17'd24215: data = 8'h1e;
      17'd24216: data = 8'h1e;
      17'd24217: data = 8'h1e;
      17'd24218: data = 8'h1a;
      17'd24219: data = 8'h13;
      17'd24220: data = 8'h0e;
      17'd24221: data = 8'h0a;
      17'd24222: data = 8'h02;
      17'd24223: data = 8'hfc;
      17'd24224: data = 8'hfd;
      17'd24225: data = 8'hfc;
      17'd24226: data = 8'hf5;
      17'd24227: data = 8'hf2;
      17'd24228: data = 8'hf2;
      17'd24229: data = 8'hed;
      17'd24230: data = 8'he7;
      17'd24231: data = 8'he9;
      17'd24232: data = 8'hec;
      17'd24233: data = 8'heb;
      17'd24234: data = 8'he7;
      17'd24235: data = 8'he9;
      17'd24236: data = 8'he7;
      17'd24237: data = 8'he7;
      17'd24238: data = 8'heb;
      17'd24239: data = 8'hf1;
      17'd24240: data = 8'hf4;
      17'd24241: data = 8'hf2;
      17'd24242: data = 8'hf6;
      17'd24243: data = 8'hfa;
      17'd24244: data = 8'hf4;
      17'd24245: data = 8'hf1;
      17'd24246: data = 8'hf4;
      17'd24247: data = 8'hf4;
      17'd24248: data = 8'hef;
      17'd24249: data = 8'hf2;
      17'd24250: data = 8'hf4;
      17'd24251: data = 8'hf1;
      17'd24252: data = 8'hf2;
      17'd24253: data = 8'hf6;
      17'd24254: data = 8'hf5;
      17'd24255: data = 8'hf6;
      17'd24256: data = 8'hfd;
      17'd24257: data = 8'h02;
      17'd24258: data = 8'h06;
      17'd24259: data = 8'h0d;
      17'd24260: data = 8'h15;
      17'd24261: data = 8'h1a;
      17'd24262: data = 8'h1f;
      17'd24263: data = 8'h24;
      17'd24264: data = 8'h27;
      17'd24265: data = 8'h24;
      17'd24266: data = 8'h24;
      17'd24267: data = 8'h24;
      17'd24268: data = 8'h1f;
      17'd24269: data = 8'h1c;
      17'd24270: data = 8'h1b;
      17'd24271: data = 8'h19;
      17'd24272: data = 8'h13;
      17'd24273: data = 8'h0d;
      17'd24274: data = 8'h0c;
      17'd24275: data = 8'h06;
      17'd24276: data = 8'h04;
      17'd24277: data = 8'h04;
      17'd24278: data = 8'h00;
      17'd24279: data = 8'hfd;
      17'd24280: data = 8'hfd;
      17'd24281: data = 8'hfa;
      17'd24282: data = 8'hf6;
      17'd24283: data = 8'hfa;
      17'd24284: data = 8'hfa;
      17'd24285: data = 8'hf6;
      17'd24286: data = 8'hf6;
      17'd24287: data = 8'hf9;
      17'd24288: data = 8'hf9;
      17'd24289: data = 8'hfc;
      17'd24290: data = 8'hfd;
      17'd24291: data = 8'hfd;
      17'd24292: data = 8'hfe;
      17'd24293: data = 8'hfe;
      17'd24294: data = 8'hfe;
      17'd24295: data = 8'hfd;
      17'd24296: data = 8'hfe;
      17'd24297: data = 8'hfe;
      17'd24298: data = 8'h01;
      17'd24299: data = 8'h00;
      17'd24300: data = 8'h00;
      17'd24301: data = 8'h01;
      17'd24302: data = 8'h01;
      17'd24303: data = 8'h01;
      17'd24304: data = 8'h02;
      17'd24305: data = 8'h02;
      17'd24306: data = 8'h01;
      17'd24307: data = 8'h02;
      17'd24308: data = 8'h02;
      17'd24309: data = 8'h02;
      17'd24310: data = 8'h04;
      17'd24311: data = 8'h05;
      17'd24312: data = 8'h0c;
      17'd24313: data = 8'h0e;
      17'd24314: data = 8'h11;
      17'd24315: data = 8'h04;
      17'd24316: data = 8'h01;
      17'd24317: data = 8'h0d;
      17'd24318: data = 8'h0c;
      17'd24319: data = 8'h06;
      17'd24320: data = 8'h11;
      17'd24321: data = 8'h0d;
      17'd24322: data = 8'h02;
      17'd24323: data = 8'h06;
      17'd24324: data = 8'h04;
      17'd24325: data = 8'hf4;
      17'd24326: data = 8'hf2;
      17'd24327: data = 8'hf9;
      17'd24328: data = 8'hf6;
      17'd24329: data = 8'hec;
      17'd24330: data = 8'hec;
      17'd24331: data = 8'hf4;
      17'd24332: data = 8'hef;
      17'd24333: data = 8'he4;
      17'd24334: data = 8'he4;
      17'd24335: data = 8'he5;
      17'd24336: data = 8'hde;
      17'd24337: data = 8'he3;
      17'd24338: data = 8'hef;
      17'd24339: data = 8'hec;
      17'd24340: data = 8'he4;
      17'd24341: data = 8'he9;
      17'd24342: data = 8'he9;
      17'd24343: data = 8'he4;
      17'd24344: data = 8'he5;
      17'd24345: data = 8'he5;
      17'd24346: data = 8'he7;
      17'd24347: data = 8'hec;
      17'd24348: data = 8'hed;
      17'd24349: data = 8'heb;
      17'd24350: data = 8'hef;
      17'd24351: data = 8'hef;
      17'd24352: data = 8'he7;
      17'd24353: data = 8'heb;
      17'd24354: data = 8'hf4;
      17'd24355: data = 8'hf4;
      17'd24356: data = 8'hef;
      17'd24357: data = 8'hf4;
      17'd24358: data = 8'hf9;
      17'd24359: data = 8'hf5;
      17'd24360: data = 8'hf4;
      17'd24361: data = 8'hf9;
      17'd24362: data = 8'hf9;
      17'd24363: data = 8'hf2;
      17'd24364: data = 8'hf4;
      17'd24365: data = 8'hfc;
      17'd24366: data = 8'hf4;
      17'd24367: data = 8'hf1;
      17'd24368: data = 8'hf6;
      17'd24369: data = 8'hfc;
      17'd24370: data = 8'hf6;
      17'd24371: data = 8'hf6;
      17'd24372: data = 8'hfe;
      17'd24373: data = 8'h05;
      17'd24374: data = 8'h06;
      17'd24375: data = 8'h0a;
      17'd24376: data = 8'h0a;
      17'd24377: data = 8'h05;
      17'd24378: data = 8'h06;
      17'd24379: data = 8'h09;
      17'd24380: data = 8'h05;
      17'd24381: data = 8'h02;
      17'd24382: data = 8'h01;
      17'd24383: data = 8'h00;
      17'd24384: data = 8'hfe;
      17'd24385: data = 8'h00;
      17'd24386: data = 8'h02;
      17'd24387: data = 8'h00;
      17'd24388: data = 8'hfe;
      17'd24389: data = 8'h00;
      17'd24390: data = 8'hfe;
      17'd24391: data = 8'hfe;
      17'd24392: data = 8'h01;
      17'd24393: data = 8'h04;
      17'd24394: data = 8'h02;
      17'd24395: data = 8'h02;
      17'd24396: data = 8'h04;
      17'd24397: data = 8'h05;
      17'd24398: data = 8'h09;
      17'd24399: data = 8'h09;
      17'd24400: data = 8'h09;
      17'd24401: data = 8'h09;
      17'd24402: data = 8'h06;
      17'd24403: data = 8'h06;
      17'd24404: data = 8'h0a;
      17'd24405: data = 8'h0a;
      17'd24406: data = 8'h09;
      17'd24407: data = 8'h0e;
      17'd24408: data = 8'h0e;
      17'd24409: data = 8'h0a;
      17'd24410: data = 8'h0a;
      17'd24411: data = 8'h0a;
      17'd24412: data = 8'h06;
      17'd24413: data = 8'h09;
      17'd24414: data = 8'h0c;
      17'd24415: data = 8'h06;
      17'd24416: data = 8'h05;
      17'd24417: data = 8'h05;
      17'd24418: data = 8'h04;
      17'd24419: data = 8'h04;
      17'd24420: data = 8'h06;
      17'd24421: data = 8'h09;
      17'd24422: data = 8'h09;
      17'd24423: data = 8'h0c;
      17'd24424: data = 8'h11;
      17'd24425: data = 8'h0c;
      17'd24426: data = 8'h02;
      17'd24427: data = 8'h01;
      17'd24428: data = 8'h01;
      17'd24429: data = 8'hf9;
      17'd24430: data = 8'hfa;
      17'd24431: data = 8'hfd;
      17'd24432: data = 8'hf2;
      17'd24433: data = 8'hec;
      17'd24434: data = 8'hf6;
      17'd24435: data = 8'hf9;
      17'd24436: data = 8'hed;
      17'd24437: data = 8'hf6;
      17'd24438: data = 8'h02;
      17'd24439: data = 8'hfe;
      17'd24440: data = 8'hfd;
      17'd24441: data = 8'h06;
      17'd24442: data = 8'h0e;
      17'd24443: data = 8'h0c;
      17'd24444: data = 8'h12;
      17'd24445: data = 8'h1c;
      17'd24446: data = 8'h1f;
      17'd24447: data = 8'h1e;
      17'd24448: data = 8'h22;
      17'd24449: data = 8'h26;
      17'd24450: data = 8'h1f;
      17'd24451: data = 8'h1e;
      17'd24452: data = 8'h1b;
      17'd24453: data = 8'h13;
      17'd24454: data = 8'h0c;
      17'd24455: data = 8'h05;
      17'd24456: data = 8'h01;
      17'd24457: data = 8'hfd;
      17'd24458: data = 8'hfc;
      17'd24459: data = 8'hf6;
      17'd24460: data = 8'hf2;
      17'd24461: data = 8'hf5;
      17'd24462: data = 8'hf5;
      17'd24463: data = 8'hed;
      17'd24464: data = 8'hec;
      17'd24465: data = 8'hf2;
      17'd24466: data = 8'hef;
      17'd24467: data = 8'hec;
      17'd24468: data = 8'hf2;
      17'd24469: data = 8'hf4;
      17'd24470: data = 8'hef;
      17'd24471: data = 8'hf1;
      17'd24472: data = 8'hf5;
      17'd24473: data = 8'hf2;
      17'd24474: data = 8'hed;
      17'd24475: data = 8'hf1;
      17'd24476: data = 8'hf2;
      17'd24477: data = 8'hec;
      17'd24478: data = 8'he9;
      17'd24479: data = 8'heb;
      17'd24480: data = 8'hec;
      17'd24481: data = 8'heb;
      17'd24482: data = 8'hec;
      17'd24483: data = 8'hef;
      17'd24484: data = 8'hef;
      17'd24485: data = 8'hf1;
      17'd24486: data = 8'hf4;
      17'd24487: data = 8'hf5;
      17'd24488: data = 8'hf9;
      17'd24489: data = 8'hfd;
      17'd24490: data = 8'h04;
      17'd24491: data = 8'h05;
      17'd24492: data = 8'h0a;
      17'd24493: data = 8'h11;
      17'd24494: data = 8'h13;
      17'd24495: data = 8'h16;
      17'd24496: data = 8'h1b;
      17'd24497: data = 8'h1e;
      17'd24498: data = 8'h1e;
      17'd24499: data = 8'h1f;
      17'd24500: data = 8'h1e;
      17'd24501: data = 8'h1f;
      17'd24502: data = 8'h1c;
      17'd24503: data = 8'h1a;
      17'd24504: data = 8'h19;
      17'd24505: data = 8'h15;
      17'd24506: data = 8'h12;
      17'd24507: data = 8'h0e;
      17'd24508: data = 8'h0c;
      17'd24509: data = 8'h0a;
      17'd24510: data = 8'h06;
      17'd24511: data = 8'h04;
      17'd24512: data = 8'h04;
      17'd24513: data = 8'h04;
      17'd24514: data = 8'h01;
      17'd24515: data = 8'h01;
      17'd24516: data = 8'h01;
      17'd24517: data = 8'h01;
      17'd24518: data = 8'h01;
      17'd24519: data = 8'h00;
      17'd24520: data = 8'h01;
      17'd24521: data = 8'h00;
      17'd24522: data = 8'h00;
      17'd24523: data = 8'h01;
      17'd24524: data = 8'h02;
      17'd24525: data = 8'h02;
      17'd24526: data = 8'h00;
      17'd24527: data = 8'h01;
      17'd24528: data = 8'h01;
      17'd24529: data = 8'h00;
      17'd24530: data = 8'h00;
      17'd24531: data = 8'hfe;
      17'd24532: data = 8'h00;
      17'd24533: data = 8'hfe;
      17'd24534: data = 8'hfc;
      17'd24535: data = 8'hfc;
      17'd24536: data = 8'hfa;
      17'd24537: data = 8'hfc;
      17'd24538: data = 8'hf9;
      17'd24539: data = 8'hfa;
      17'd24540: data = 8'hfc;
      17'd24541: data = 8'hfe;
      17'd24542: data = 8'h00;
      17'd24543: data = 8'h02;
      17'd24544: data = 8'h05;
      17'd24545: data = 8'h09;
      17'd24546: data = 8'h0a;
      17'd24547: data = 8'h09;
      17'd24548: data = 8'h09;
      17'd24549: data = 8'h0a;
      17'd24550: data = 8'h09;
      17'd24551: data = 8'h0a;
      17'd24552: data = 8'h0a;
      17'd24553: data = 8'h06;
      17'd24554: data = 8'h05;
      17'd24555: data = 8'h00;
      17'd24556: data = 8'h00;
      17'd24557: data = 8'hfd;
      17'd24558: data = 8'hfa;
      17'd24559: data = 8'hf6;
      17'd24560: data = 8'hf5;
      17'd24561: data = 8'hf6;
      17'd24562: data = 8'hf4;
      17'd24563: data = 8'hf4;
      17'd24564: data = 8'hf2;
      17'd24565: data = 8'hf1;
      17'd24566: data = 8'hef;
      17'd24567: data = 8'hef;
      17'd24568: data = 8'hf1;
      17'd24569: data = 8'hef;
      17'd24570: data = 8'hf2;
      17'd24571: data = 8'hf1;
      17'd24572: data = 8'hef;
      17'd24573: data = 8'hef;
      17'd24574: data = 8'hed;
      17'd24575: data = 8'hed;
      17'd24576: data = 8'hec;
      17'd24577: data = 8'heb;
      17'd24578: data = 8'heb;
      17'd24579: data = 8'he9;
      17'd24580: data = 8'he5;
      17'd24581: data = 8'he4;
      17'd24582: data = 8'he4;
      17'd24583: data = 8'he3;
      17'd24584: data = 8'he2;
      17'd24585: data = 8'he2;
      17'd24586: data = 8'he3;
      17'd24587: data = 8'he3;
      17'd24588: data = 8'he3;
      17'd24589: data = 8'he5;
      17'd24590: data = 8'he7;
      17'd24591: data = 8'he9;
      17'd24592: data = 8'hec;
      17'd24593: data = 8'hec;
      17'd24594: data = 8'hed;
      17'd24595: data = 8'hef;
      17'd24596: data = 8'hf1;
      17'd24597: data = 8'hf1;
      17'd24598: data = 8'hf1;
      17'd24599: data = 8'hf2;
      17'd24600: data = 8'hf4;
      17'd24601: data = 8'hf5;
      17'd24602: data = 8'hf5;
      17'd24603: data = 8'hfa;
      17'd24604: data = 8'hfc;
      17'd24605: data = 8'hfc;
      17'd24606: data = 8'h00;
      17'd24607: data = 8'h00;
      17'd24608: data = 8'h01;
      17'd24609: data = 8'h04;
      17'd24610: data = 8'h05;
      17'd24611: data = 8'h09;
      17'd24612: data = 8'h0a;
      17'd24613: data = 8'h0c;
      17'd24614: data = 8'h0c;
      17'd24615: data = 8'h0c;
      17'd24616: data = 8'h0d;
      17'd24617: data = 8'h0d;
      17'd24618: data = 8'h0d;
      17'd24619: data = 8'h0c;
      17'd24620: data = 8'h0a;
      17'd24621: data = 8'h06;
      17'd24622: data = 8'h05;
      17'd24623: data = 8'h06;
      17'd24624: data = 8'h06;
      17'd24625: data = 8'h09;
      17'd24626: data = 8'h06;
      17'd24627: data = 8'h06;
      17'd24628: data = 8'h0a;
      17'd24629: data = 8'h0a;
      17'd24630: data = 8'h05;
      17'd24631: data = 8'h09;
      17'd24632: data = 8'h09;
      17'd24633: data = 8'h06;
      17'd24634: data = 8'h06;
      17'd24635: data = 8'h04;
      17'd24636: data = 8'h02;
      17'd24637: data = 8'h04;
      17'd24638: data = 8'h05;
      17'd24639: data = 8'h02;
      17'd24640: data = 8'h06;
      17'd24641: data = 8'h09;
      17'd24642: data = 8'h04;
      17'd24643: data = 8'h04;
      17'd24644: data = 8'h04;
      17'd24645: data = 8'h04;
      17'd24646: data = 8'h04;
      17'd24647: data = 8'h04;
      17'd24648: data = 8'h04;
      17'd24649: data = 8'h06;
      17'd24650: data = 8'h01;
      17'd24651: data = 8'h00;
      17'd24652: data = 8'h04;
      17'd24653: data = 8'h00;
      17'd24654: data = 8'h00;
      17'd24655: data = 8'h05;
      17'd24656: data = 8'h0a;
      17'd24657: data = 8'h04;
      17'd24658: data = 8'h05;
      17'd24659: data = 8'h0c;
      17'd24660: data = 8'h0a;
      17'd24661: data = 8'h04;
      17'd24662: data = 8'h05;
      17'd24663: data = 8'h05;
      17'd24664: data = 8'h01;
      17'd24665: data = 8'h04;
      17'd24666: data = 8'h02;
      17'd24667: data = 8'h00;
      17'd24668: data = 8'hfc;
      17'd24669: data = 8'hf6;
      17'd24670: data = 8'hf5;
      17'd24671: data = 8'hf5;
      17'd24672: data = 8'hf6;
      17'd24673: data = 8'hfa;
      17'd24674: data = 8'hfe;
      17'd24675: data = 8'h02;
      17'd24676: data = 8'h09;
      17'd24677: data = 8'h0c;
      17'd24678: data = 8'h0a;
      17'd24679: data = 8'h0e;
      17'd24680: data = 8'h16;
      17'd24681: data = 8'h16;
      17'd24682: data = 8'h16;
      17'd24683: data = 8'h1b;
      17'd24684: data = 8'h15;
      17'd24685: data = 8'h0e;
      17'd24686: data = 8'h12;
      17'd24687: data = 8'h0e;
      17'd24688: data = 8'h09;
      17'd24689: data = 8'h06;
      17'd24690: data = 8'h05;
      17'd24691: data = 8'h01;
      17'd24692: data = 8'hfd;
      17'd24693: data = 8'hf9;
      17'd24694: data = 8'hf2;
      17'd24695: data = 8'hf1;
      17'd24696: data = 8'hf1;
      17'd24697: data = 8'hed;
      17'd24698: data = 8'hec;
      17'd24699: data = 8'hec;
      17'd24700: data = 8'hef;
      17'd24701: data = 8'hef;
      17'd24702: data = 8'hf4;
      17'd24703: data = 8'hf6;
      17'd24704: data = 8'hf9;
      17'd24705: data = 8'hf9;
      17'd24706: data = 8'hfa;
      17'd24707: data = 8'hfc;
      17'd24708: data = 8'hf9;
      17'd24709: data = 8'hf5;
      17'd24710: data = 8'hf4;
      17'd24711: data = 8'hf5;
      17'd24712: data = 8'hf2;
      17'd24713: data = 8'hf1;
      17'd24714: data = 8'hf1;
      17'd24715: data = 8'hef;
      17'd24716: data = 8'hef;
      17'd24717: data = 8'hf4;
      17'd24718: data = 8'hf6;
      17'd24719: data = 8'hf5;
      17'd24720: data = 8'hf5;
      17'd24721: data = 8'hf5;
      17'd24722: data = 8'hf6;
      17'd24723: data = 8'hfa;
      17'd24724: data = 8'hfa;
      17'd24725: data = 8'hfd;
      17'd24726: data = 8'h01;
      17'd24727: data = 8'h04;
      17'd24728: data = 8'h09;
      17'd24729: data = 8'h0d;
      17'd24730: data = 8'h11;
      17'd24731: data = 8'h15;
      17'd24732: data = 8'h1a;
      17'd24733: data = 8'h1c;
      17'd24734: data = 8'h1b;
      17'd24735: data = 8'h1b;
      17'd24736: data = 8'h1b;
      17'd24737: data = 8'h16;
      17'd24738: data = 8'h15;
      17'd24739: data = 8'h13;
      17'd24740: data = 8'h0e;
      17'd24741: data = 8'h0d;
      17'd24742: data = 8'h09;
      17'd24743: data = 8'h09;
      17'd24744: data = 8'h05;
      17'd24745: data = 8'h02;
      17'd24746: data = 8'h01;
      17'd24747: data = 8'h02;
      17'd24748: data = 8'h05;
      17'd24749: data = 8'h06;
      17'd24750: data = 8'h09;
      17'd24751: data = 8'h0a;
      17'd24752: data = 8'h0c;
      17'd24753: data = 8'h09;
      17'd24754: data = 8'h09;
      17'd24755: data = 8'h0a;
      17'd24756: data = 8'h09;
      17'd24757: data = 8'h09;
      17'd24758: data = 8'h0a;
      17'd24759: data = 8'h0a;
      17'd24760: data = 8'h09;
      17'd24761: data = 8'h06;
      17'd24762: data = 8'h05;
      17'd24763: data = 8'h02;
      17'd24764: data = 8'h01;
      17'd24765: data = 8'hfe;
      17'd24766: data = 8'hfd;
      17'd24767: data = 8'hfa;
      17'd24768: data = 8'hfa;
      17'd24769: data = 8'hf9;
      17'd24770: data = 8'hf9;
      17'd24771: data = 8'hf9;
      17'd24772: data = 8'hf9;
      17'd24773: data = 8'hfa;
      17'd24774: data = 8'hfd;
      17'd24775: data = 8'h00;
      17'd24776: data = 8'h01;
      17'd24777: data = 8'h02;
      17'd24778: data = 8'h02;
      17'd24779: data = 8'h01;
      17'd24780: data = 8'h00;
      17'd24781: data = 8'h01;
      17'd24782: data = 8'h01;
      17'd24783: data = 8'h01;
      17'd24784: data = 8'h02;
      17'd24785: data = 8'h01;
      17'd24786: data = 8'hfe;
      17'd24787: data = 8'h01;
      17'd24788: data = 8'h01;
      17'd24789: data = 8'hfe;
      17'd24790: data = 8'hfa;
      17'd24791: data = 8'hfc;
      17'd24792: data = 8'hfc;
      17'd24793: data = 8'hf9;
      17'd24794: data = 8'hfa;
      17'd24795: data = 8'hfa;
      17'd24796: data = 8'hf6;
      17'd24797: data = 8'hf5;
      17'd24798: data = 8'hf6;
      17'd24799: data = 8'hf5;
      17'd24800: data = 8'hf4;
      17'd24801: data = 8'hf2;
      17'd24802: data = 8'hf2;
      17'd24803: data = 8'hf4;
      17'd24804: data = 8'hf2;
      17'd24805: data = 8'hf2;
      17'd24806: data = 8'hf2;
      17'd24807: data = 8'hef;
      17'd24808: data = 8'hec;
      17'd24809: data = 8'heb;
      17'd24810: data = 8'he9;
      17'd24811: data = 8'he5;
      17'd24812: data = 8'he3;
      17'd24813: data = 8'he4;
      17'd24814: data = 8'he4;
      17'd24815: data = 8'he3;
      17'd24816: data = 8'he0;
      17'd24817: data = 8'he0;
      17'd24818: data = 8'he3;
      17'd24819: data = 8'he3;
      17'd24820: data = 8'he4;
      17'd24821: data = 8'he4;
      17'd24822: data = 8'he4;
      17'd24823: data = 8'he4;
      17'd24824: data = 8'he5;
      17'd24825: data = 8'he7;
      17'd24826: data = 8'he9;
      17'd24827: data = 8'he9;
      17'd24828: data = 8'heb;
      17'd24829: data = 8'hef;
      17'd24830: data = 8'hef;
      17'd24831: data = 8'hf2;
      17'd24832: data = 8'hf2;
      17'd24833: data = 8'hf4;
      17'd24834: data = 8'hf5;
      17'd24835: data = 8'hf6;
      17'd24836: data = 8'hf9;
      17'd24837: data = 8'hf9;
      17'd24838: data = 8'hfa;
      17'd24839: data = 8'hfa;
      17'd24840: data = 8'hfc;
      17'd24841: data = 8'hfc;
      17'd24842: data = 8'h00;
      17'd24843: data = 8'h02;
      17'd24844: data = 8'h05;
      17'd24845: data = 8'h05;
      17'd24846: data = 8'h09;
      17'd24847: data = 8'h0d;
      17'd24848: data = 8'h0d;
      17'd24849: data = 8'h11;
      17'd24850: data = 8'h11;
      17'd24851: data = 8'h0e;
      17'd24852: data = 8'h0c;
      17'd24853: data = 8'h0a;
      17'd24854: data = 8'h09;
      17'd24855: data = 8'h05;
      17'd24856: data = 8'h06;
      17'd24857: data = 8'h06;
      17'd24858: data = 8'h0a;
      17'd24859: data = 8'h09;
      17'd24860: data = 8'h06;
      17'd24861: data = 8'h0a;
      17'd24862: data = 8'h06;
      17'd24863: data = 8'h02;
      17'd24864: data = 8'h02;
      17'd24865: data = 8'h04;
      17'd24866: data = 8'h06;
      17'd24867: data = 8'h06;
      17'd24868: data = 8'h09;
      17'd24869: data = 8'h09;
      17'd24870: data = 8'h0c;
      17'd24871: data = 8'h0d;
      17'd24872: data = 8'h0d;
      17'd24873: data = 8'h04;
      17'd24874: data = 8'hfa;
      17'd24875: data = 8'h0a;
      17'd24876: data = 8'h16;
      17'd24877: data = 8'h0a;
      17'd24878: data = 8'hfe;
      17'd24879: data = 8'h02;
      17'd24880: data = 8'h06;
      17'd24881: data = 8'h0a;
      17'd24882: data = 8'h09;
      17'd24883: data = 8'h00;
      17'd24884: data = 8'h06;
      17'd24885: data = 8'h13;
      17'd24886: data = 8'h0a;
      17'd24887: data = 8'h06;
      17'd24888: data = 8'h0d;
      17'd24889: data = 8'h11;
      17'd24890: data = 8'h0d;
      17'd24891: data = 8'h0c;
      17'd24892: data = 8'h0d;
      17'd24893: data = 8'h0c;
      17'd24894: data = 8'h0a;
      17'd24895: data = 8'h09;
      17'd24896: data = 8'h0a;
      17'd24897: data = 8'h0c;
      17'd24898: data = 8'h0a;
      17'd24899: data = 8'h05;
      17'd24900: data = 8'h06;
      17'd24901: data = 8'h05;
      17'd24902: data = 8'hfd;
      17'd24903: data = 8'hfa;
      17'd24904: data = 8'hfc;
      17'd24905: data = 8'hfd;
      17'd24906: data = 8'hfa;
      17'd24907: data = 8'hf5;
      17'd24908: data = 8'hf4;
      17'd24909: data = 8'hf6;
      17'd24910: data = 8'hfa;
      17'd24911: data = 8'h00;
      17'd24912: data = 8'h02;
      17'd24913: data = 8'h02;
      17'd24914: data = 8'h05;
      17'd24915: data = 8'h04;
      17'd24916: data = 8'h02;
      17'd24917: data = 8'h05;
      17'd24918: data = 8'h06;
      17'd24919: data = 8'h06;
      17'd24920: data = 8'h0c;
      17'd24921: data = 8'h0d;
      17'd24922: data = 8'h05;
      17'd24923: data = 8'h05;
      17'd24924: data = 8'h06;
      17'd24925: data = 8'h02;
      17'd24926: data = 8'h00;
      17'd24927: data = 8'h05;
      17'd24928: data = 8'h0a;
      17'd24929: data = 8'h0a;
      17'd24930: data = 8'h06;
      17'd24931: data = 8'h04;
      17'd24932: data = 8'h06;
      17'd24933: data = 8'h06;
      17'd24934: data = 8'h04;
      17'd24935: data = 8'h06;
      17'd24936: data = 8'h0a;
      17'd24937: data = 8'h0a;
      17'd24938: data = 8'h0a;
      17'd24939: data = 8'h0d;
      17'd24940: data = 8'h0d;
      17'd24941: data = 8'h0c;
      17'd24942: data = 8'h0c;
      17'd24943: data = 8'h0a;
      17'd24944: data = 8'h0a;
      17'd24945: data = 8'h06;
      17'd24946: data = 8'h04;
      17'd24947: data = 8'h01;
      17'd24948: data = 8'h00;
      17'd24949: data = 8'hfc;
      17'd24950: data = 8'hfa;
      17'd24951: data = 8'hf9;
      17'd24952: data = 8'hf6;
      17'd24953: data = 8'hf5;
      17'd24954: data = 8'hf6;
      17'd24955: data = 8'hf6;
      17'd24956: data = 8'hf4;
      17'd24957: data = 8'hf2;
      17'd24958: data = 8'hf2;
      17'd24959: data = 8'hf2;
      17'd24960: data = 8'hf1;
      17'd24961: data = 8'hf1;
      17'd24962: data = 8'hf1;
      17'd24963: data = 8'hf1;
      17'd24964: data = 8'hf4;
      17'd24965: data = 8'hf4;
      17'd24966: data = 8'hf4;
      17'd24967: data = 8'hfa;
      17'd24968: data = 8'hfd;
      17'd24969: data = 8'hfd;
      17'd24970: data = 8'h02;
      17'd24971: data = 8'h02;
      17'd24972: data = 8'h04;
      17'd24973: data = 8'h04;
      17'd24974: data = 8'h02;
      17'd24975: data = 8'h02;
      17'd24976: data = 8'h01;
      17'd24977: data = 8'hfe;
      17'd24978: data = 8'hfe;
      17'd24979: data = 8'h01;
      17'd24980: data = 8'h01;
      17'd24981: data = 8'h02;
      17'd24982: data = 8'h06;
      17'd24983: data = 8'h09;
      17'd24984: data = 8'h0a;
      17'd24985: data = 8'h0d;
      17'd24986: data = 8'h0d;
      17'd24987: data = 8'h0e;
      17'd24988: data = 8'h13;
      17'd24989: data = 8'h13;
      17'd24990: data = 8'h12;
      17'd24991: data = 8'h13;
      17'd24992: data = 8'h13;
      17'd24993: data = 8'h12;
      17'd24994: data = 8'h11;
      17'd24995: data = 8'h11;
      17'd24996: data = 8'h0d;
      17'd24997: data = 8'h0d;
      17'd24998: data = 8'h0d;
      17'd24999: data = 8'h0c;
      17'd25000: data = 8'h0c;
      17'd25001: data = 8'h09;
      17'd25002: data = 8'h05;
      17'd25003: data = 8'h04;
      17'd25004: data = 8'h02;
      17'd25005: data = 8'h01;
      17'd25006: data = 8'h00;
      17'd25007: data = 8'hfd;
      17'd25008: data = 8'hfc;
      17'd25009: data = 8'hfd;
      17'd25010: data = 8'hfe;
      17'd25011: data = 8'hfa;
      17'd25012: data = 8'hfa;
      17'd25013: data = 8'hfa;
      17'd25014: data = 8'hfc;
      17'd25015: data = 8'hfd;
      17'd25016: data = 8'hf9;
      17'd25017: data = 8'hf9;
      17'd25018: data = 8'hf9;
      17'd25019: data = 8'hf6;
      17'd25020: data = 8'hf6;
      17'd25021: data = 8'hf4;
      17'd25022: data = 8'hf5;
      17'd25023: data = 8'hf4;
      17'd25024: data = 8'hf4;
      17'd25025: data = 8'hf9;
      17'd25026: data = 8'hf9;
      17'd25027: data = 8'hf9;
      17'd25028: data = 8'hfd;
      17'd25029: data = 8'h00;
      17'd25030: data = 8'hfe;
      17'd25031: data = 8'hfc;
      17'd25032: data = 8'hfd;
      17'd25033: data = 8'hfc;
      17'd25034: data = 8'hf9;
      17'd25035: data = 8'hf6;
      17'd25036: data = 8'hf9;
      17'd25037: data = 8'hf6;
      17'd25038: data = 8'hf5;
      17'd25039: data = 8'hf4;
      17'd25040: data = 8'hf5;
      17'd25041: data = 8'hf6;
      17'd25042: data = 8'hf6;
      17'd25043: data = 8'hf5;
      17'd25044: data = 8'hf5;
      17'd25045: data = 8'hf4;
      17'd25046: data = 8'hf1;
      17'd25047: data = 8'hef;
      17'd25048: data = 8'hec;
      17'd25049: data = 8'hec;
      17'd25050: data = 8'heb;
      17'd25051: data = 8'he9;
      17'd25052: data = 8'he9;
      17'd25053: data = 8'hec;
      17'd25054: data = 8'heb;
      17'd25055: data = 8'hec;
      17'd25056: data = 8'heb;
      17'd25057: data = 8'he9;
      17'd25058: data = 8'heb;
      17'd25059: data = 8'he9;
      17'd25060: data = 8'he9;
      17'd25061: data = 8'he7;
      17'd25062: data = 8'he4;
      17'd25063: data = 8'he4;
      17'd25064: data = 8'he4;
      17'd25065: data = 8'he3;
      17'd25066: data = 8'he3;
      17'd25067: data = 8'he2;
      17'd25068: data = 8'he3;
      17'd25069: data = 8'he5;
      17'd25070: data = 8'he9;
      17'd25071: data = 8'he9;
      17'd25072: data = 8'he9;
      17'd25073: data = 8'heb;
      17'd25074: data = 8'heb;
      17'd25075: data = 8'hed;
      17'd25076: data = 8'hef;
      17'd25077: data = 8'hf1;
      17'd25078: data = 8'hf2;
      17'd25079: data = 8'hf1;
      17'd25080: data = 8'hf4;
      17'd25081: data = 8'hf5;
      17'd25082: data = 8'hf5;
      17'd25083: data = 8'hf9;
      17'd25084: data = 8'hfa;
      17'd25085: data = 8'hfc;
      17'd25086: data = 8'hfd;
      17'd25087: data = 8'h00;
      17'd25088: data = 8'h00;
      17'd25089: data = 8'hfe;
      17'd25090: data = 8'h00;
      17'd25091: data = 8'h02;
      17'd25092: data = 8'h04;
      17'd25093: data = 8'h06;
      17'd25094: data = 8'h0a;
      17'd25095: data = 8'h0a;
      17'd25096: data = 8'h0a;
      17'd25097: data = 8'h0d;
      17'd25098: data = 8'h0e;
      17'd25099: data = 8'h12;
      17'd25100: data = 8'h12;
      17'd25101: data = 8'h15;
      17'd25102: data = 8'h16;
      17'd25103: data = 8'h16;
      17'd25104: data = 8'h15;
      17'd25105: data = 8'h15;
      17'd25106: data = 8'h12;
      17'd25107: data = 8'h0e;
      17'd25108: data = 8'h12;
      17'd25109: data = 8'h11;
      17'd25110: data = 8'h0e;
      17'd25111: data = 8'h0d;
      17'd25112: data = 8'h0e;
      17'd25113: data = 8'h11;
      17'd25114: data = 8'h0e;
      17'd25115: data = 8'h11;
      17'd25116: data = 8'h11;
      17'd25117: data = 8'h11;
      17'd25118: data = 8'h11;
      17'd25119: data = 8'h0e;
      17'd25120: data = 8'h11;
      17'd25121: data = 8'h11;
      17'd25122: data = 8'h09;
      17'd25123: data = 8'h09;
      17'd25124: data = 8'h09;
      17'd25125: data = 8'h04;
      17'd25126: data = 8'h01;
      17'd25127: data = 8'h02;
      17'd25128: data = 8'h04;
      17'd25129: data = 8'h02;
      17'd25130: data = 8'h04;
      17'd25131: data = 8'h02;
      17'd25132: data = 8'h01;
      17'd25133: data = 8'h00;
      17'd25134: data = 8'hfd;
      17'd25135: data = 8'hfc;
      17'd25136: data = 8'hfd;
      17'd25137: data = 8'hfc;
      17'd25138: data = 8'hfe;
      17'd25139: data = 8'hfc;
      17'd25140: data = 8'hfc;
      17'd25141: data = 8'hfa;
      17'd25142: data = 8'hf5;
      17'd25143: data = 8'hf5;
      17'd25144: data = 8'hf9;
      17'd25145: data = 8'hfa;
      17'd25146: data = 8'hfd;
      17'd25147: data = 8'h00;
      17'd25148: data = 8'h04;
      17'd25149: data = 8'h05;
      17'd25150: data = 8'h01;
      17'd25151: data = 8'h00;
      17'd25152: data = 8'h09;
      17'd25153: data = 8'h0e;
      17'd25154: data = 8'h0e;
      17'd25155: data = 8'h13;
      17'd25156: data = 8'h19;
      17'd25157: data = 8'h16;
      17'd25158: data = 8'h11;
      17'd25159: data = 8'h0a;
      17'd25160: data = 8'h0a;
      17'd25161: data = 8'h0c;
      17'd25162: data = 8'h06;
      17'd25163: data = 8'h05;
      17'd25164: data = 8'h0c;
      17'd25165: data = 8'h0c;
      17'd25166: data = 8'h05;
      17'd25167: data = 8'h06;
      17'd25168: data = 8'h0a;
      17'd25169: data = 8'h0a;
      17'd25170: data = 8'h0c;
      17'd25171: data = 8'h11;
      17'd25172: data = 8'h11;
      17'd25173: data = 8'h13;
      17'd25174: data = 8'h12;
      17'd25175: data = 8'h0e;
      17'd25176: data = 8'h11;
      17'd25177: data = 8'h0a;
      17'd25178: data = 8'h04;
      17'd25179: data = 8'h04;
      17'd25180: data = 8'h02;
      17'd25181: data = 8'hfc;
      17'd25182: data = 8'hf6;
      17'd25183: data = 8'hf4;
      17'd25184: data = 8'hf2;
      17'd25185: data = 8'hef;
      17'd25186: data = 8'he9;
      17'd25187: data = 8'he9;
      17'd25188: data = 8'hec;
      17'd25189: data = 8'hec;
      17'd25190: data = 8'heb;
      17'd25191: data = 8'hec;
      17'd25192: data = 8'hf1;
      17'd25193: data = 8'hef;
      17'd25194: data = 8'hef;
      17'd25195: data = 8'hf2;
      17'd25196: data = 8'hf4;
      17'd25197: data = 8'hf4;
      17'd25198: data = 8'hf4;
      17'd25199: data = 8'hf6;
      17'd25200: data = 8'hf6;
      17'd25201: data = 8'hf6;
      17'd25202: data = 8'hf5;
      17'd25203: data = 8'hf4;
      17'd25204: data = 8'hf9;
      17'd25205: data = 8'hf9;
      17'd25206: data = 8'hfa;
      17'd25207: data = 8'h00;
      17'd25208: data = 8'h01;
      17'd25209: data = 8'h02;
      17'd25210: data = 8'h06;
      17'd25211: data = 8'h0a;
      17'd25212: data = 8'h0d;
      17'd25213: data = 8'h0d;
      17'd25214: data = 8'h0a;
      17'd25215: data = 8'h0d;
      17'd25216: data = 8'h0e;
      17'd25217: data = 8'h0d;
      17'd25218: data = 8'h0c;
      17'd25219: data = 8'h0e;
      17'd25220: data = 8'h12;
      17'd25221: data = 8'h11;
      17'd25222: data = 8'h11;
      17'd25223: data = 8'h12;
      17'd25224: data = 8'h13;
      17'd25225: data = 8'h16;
      17'd25226: data = 8'h15;
      17'd25227: data = 8'h15;
      17'd25228: data = 8'h13;
      17'd25229: data = 8'h12;
      17'd25230: data = 8'h12;
      17'd25231: data = 8'h12;
      17'd25232: data = 8'h0e;
      17'd25233: data = 8'h0a;
      17'd25234: data = 8'h0a;
      17'd25235: data = 8'h06;
      17'd25236: data = 8'h06;
      17'd25237: data = 8'h04;
      17'd25238: data = 8'h02;
      17'd25239: data = 8'h01;
      17'd25240: data = 8'h00;
      17'd25241: data = 8'hfe;
      17'd25242: data = 8'hfc;
      17'd25243: data = 8'hfa;
      17'd25244: data = 8'hfa;
      17'd25245: data = 8'hfc;
      17'd25246: data = 8'hfa;
      17'd25247: data = 8'hfa;
      17'd25248: data = 8'hf6;
      17'd25249: data = 8'hf6;
      17'd25250: data = 8'hf9;
      17'd25251: data = 8'hf9;
      17'd25252: data = 8'hf4;
      17'd25253: data = 8'hf2;
      17'd25254: data = 8'hf1;
      17'd25255: data = 8'hf4;
      17'd25256: data = 8'hf4;
      17'd25257: data = 8'hed;
      17'd25258: data = 8'hec;
      17'd25259: data = 8'hf1;
      17'd25260: data = 8'hf5;
      17'd25261: data = 8'hf1;
      17'd25262: data = 8'hf4;
      17'd25263: data = 8'hfa;
      17'd25264: data = 8'hfd;
      17'd25265: data = 8'hfd;
      17'd25266: data = 8'hfa;
      17'd25267: data = 8'hfd;
      17'd25268: data = 8'hfa;
      17'd25269: data = 8'hf9;
      17'd25270: data = 8'hfd;
      17'd25271: data = 8'hfd;
      17'd25272: data = 8'hf9;
      17'd25273: data = 8'hf5;
      17'd25274: data = 8'hf9;
      17'd25275: data = 8'hf9;
      17'd25276: data = 8'hf4;
      17'd25277: data = 8'hf1;
      17'd25278: data = 8'hf2;
      17'd25279: data = 8'hf5;
      17'd25280: data = 8'hf2;
      17'd25281: data = 8'hf4;
      17'd25282: data = 8'hf5;
      17'd25283: data = 8'hf4;
      17'd25284: data = 8'hf1;
      17'd25285: data = 8'hf2;
      17'd25286: data = 8'hf4;
      17'd25287: data = 8'hef;
      17'd25288: data = 8'he9;
      17'd25289: data = 8'he9;
      17'd25290: data = 8'heb;
      17'd25291: data = 8'he7;
      17'd25292: data = 8'he4;
      17'd25293: data = 8'he3;
      17'd25294: data = 8'he5;
      17'd25295: data = 8'he7;
      17'd25296: data = 8'he5;
      17'd25297: data = 8'he5;
      17'd25298: data = 8'he5;
      17'd25299: data = 8'he7;
      17'd25300: data = 8'he5;
      17'd25301: data = 8'he4;
      17'd25302: data = 8'he5;
      17'd25303: data = 8'he7;
      17'd25304: data = 8'he7;
      17'd25305: data = 8'he7;
      17'd25306: data = 8'he5;
      17'd25307: data = 8'he5;
      17'd25308: data = 8'he7;
      17'd25309: data = 8'he5;
      17'd25310: data = 8'he7;
      17'd25311: data = 8'heb;
      17'd25312: data = 8'heb;
      17'd25313: data = 8'hec;
      17'd25314: data = 8'hef;
      17'd25315: data = 8'hf2;
      17'd25316: data = 8'hf1;
      17'd25317: data = 8'hf4;
      17'd25318: data = 8'hfc;
      17'd25319: data = 8'hfd;
      17'd25320: data = 8'h00;
      17'd25321: data = 8'h02;
      17'd25322: data = 8'h06;
      17'd25323: data = 8'h06;
      17'd25324: data = 8'h06;
      17'd25325: data = 8'h0c;
      17'd25326: data = 8'h0d;
      17'd25327: data = 8'h0d;
      17'd25328: data = 8'h0c;
      17'd25329: data = 8'h0e;
      17'd25330: data = 8'h11;
      17'd25331: data = 8'h0e;
      17'd25332: data = 8'h0c;
      17'd25333: data = 8'h0d;
      17'd25334: data = 8'h11;
      17'd25335: data = 8'h0d;
      17'd25336: data = 8'h11;
      17'd25337: data = 8'h13;
      17'd25338: data = 8'h13;
      17'd25339: data = 8'h15;
      17'd25340: data = 8'h15;
      17'd25341: data = 8'h19;
      17'd25342: data = 8'h19;
      17'd25343: data = 8'h15;
      17'd25344: data = 8'h15;
      17'd25345: data = 8'h15;
      17'd25346: data = 8'h12;
      17'd25347: data = 8'h11;
      17'd25348: data = 8'h11;
      17'd25349: data = 8'h0e;
      17'd25350: data = 8'h09;
      17'd25351: data = 8'h09;
      17'd25352: data = 8'h05;
      17'd25353: data = 8'h04;
      17'd25354: data = 8'h06;
      17'd25355: data = 8'h05;
      17'd25356: data = 8'h05;
      17'd25357: data = 8'h05;
      17'd25358: data = 8'h05;
      17'd25359: data = 8'h05;
      17'd25360: data = 8'h05;
      17'd25361: data = 8'h09;
      17'd25362: data = 8'h0a;
      17'd25363: data = 8'h06;
      17'd25364: data = 8'h04;
      17'd25365: data = 8'h02;
      17'd25366: data = 8'h01;
      17'd25367: data = 8'hfc;
      17'd25368: data = 8'hfa;
      17'd25369: data = 8'hfc;
      17'd25370: data = 8'hfd;
      17'd25371: data = 8'hfe;
      17'd25372: data = 8'hfe;
      17'd25373: data = 8'hfe;
      17'd25374: data = 8'hfe;
      17'd25375: data = 8'hfa;
      17'd25376: data = 8'hfa;
      17'd25377: data = 8'h01;
      17'd25378: data = 8'h02;
      17'd25379: data = 8'h02;
      17'd25380: data = 8'h0a;
      17'd25381: data = 8'h11;
      17'd25382: data = 8'h0e;
      17'd25383: data = 8'h09;
      17'd25384: data = 8'h09;
      17'd25385: data = 8'h0c;
      17'd25386: data = 8'h0e;
      17'd25387: data = 8'h0d;
      17'd25388: data = 8'h0e;
      17'd25389: data = 8'h12;
      17'd25390: data = 8'h11;
      17'd25391: data = 8'h0d;
      17'd25392: data = 8'h0d;
      17'd25393: data = 8'h0c;
      17'd25394: data = 8'h0a;
      17'd25395: data = 8'h0c;
      17'd25396: data = 8'h12;
      17'd25397: data = 8'h15;
      17'd25398: data = 8'h0e;
      17'd25399: data = 8'h0c;
      17'd25400: data = 8'h0d;
      17'd25401: data = 8'h0c;
      17'd25402: data = 8'h06;
      17'd25403: data = 8'h05;
      17'd25404: data = 8'h06;
      17'd25405: data = 8'h0a;
      17'd25406: data = 8'h0c;
      17'd25407: data = 8'h0c;
      17'd25408: data = 8'h0a;
      17'd25409: data = 8'h09;
      17'd25410: data = 8'h02;
      17'd25411: data = 8'h01;
      17'd25412: data = 8'h02;
      17'd25413: data = 8'hfe;
      17'd25414: data = 8'hfc;
      17'd25415: data = 8'hfd;
      17'd25416: data = 8'hfa;
      17'd25417: data = 8'hf6;
      17'd25418: data = 8'hf4;
      17'd25419: data = 8'hef;
      17'd25420: data = 8'hed;
      17'd25421: data = 8'hed;
      17'd25422: data = 8'hed;
      17'd25423: data = 8'hed;
      17'd25424: data = 8'hec;
      17'd25425: data = 8'hef;
      17'd25426: data = 8'hef;
      17'd25427: data = 8'hef;
      17'd25428: data = 8'hf1;
      17'd25429: data = 8'hf1;
      17'd25430: data = 8'hf2;
      17'd25431: data = 8'hf5;
      17'd25432: data = 8'hf9;
      17'd25433: data = 8'hf9;
      17'd25434: data = 8'hf9;
      17'd25435: data = 8'hfa;
      17'd25436: data = 8'hfa;
      17'd25437: data = 8'hfd;
      17'd25438: data = 8'h00;
      17'd25439: data = 8'hfe;
      17'd25440: data = 8'h01;
      17'd25441: data = 8'h02;
      17'd25442: data = 8'h04;
      17'd25443: data = 8'h04;
      17'd25444: data = 8'h06;
      17'd25445: data = 8'h06;
      17'd25446: data = 8'h09;
      17'd25447: data = 8'h0c;
      17'd25448: data = 8'h0c;
      17'd25449: data = 8'h0d;
      17'd25450: data = 8'h11;
      17'd25451: data = 8'h13;
      17'd25452: data = 8'h16;
      17'd25453: data = 8'h16;
      17'd25454: data = 8'h15;
      17'd25455: data = 8'h15;
      17'd25456: data = 8'h16;
      17'd25457: data = 8'h13;
      17'd25458: data = 8'h12;
      17'd25459: data = 8'h12;
      17'd25460: data = 8'h11;
      17'd25461: data = 8'h12;
      17'd25462: data = 8'h11;
      17'd25463: data = 8'h0e;
      17'd25464: data = 8'h0c;
      17'd25465: data = 8'h0e;
      17'd25466: data = 8'h0d;
      17'd25467: data = 8'h0c;
      17'd25468: data = 8'h0c;
      17'd25469: data = 8'h0a;
      17'd25470: data = 8'h0a;
      17'd25471: data = 8'h09;
      17'd25472: data = 8'h06;
      17'd25473: data = 8'h04;
      17'd25474: data = 8'h02;
      17'd25475: data = 8'h00;
      17'd25476: data = 8'hfd;
      17'd25477: data = 8'hfe;
      17'd25478: data = 8'hfd;
      17'd25479: data = 8'hf9;
      17'd25480: data = 8'hfa;
      17'd25481: data = 8'hfa;
      17'd25482: data = 8'hfa;
      17'd25483: data = 8'hfa;
      17'd25484: data = 8'hf9;
      17'd25485: data = 8'hfc;
      17'd25486: data = 8'hf6;
      17'd25487: data = 8'hf4;
      17'd25488: data = 8'hf1;
      17'd25489: data = 8'hef;
      17'd25490: data = 8'hef;
      17'd25491: data = 8'hec;
      17'd25492: data = 8'hed;
      17'd25493: data = 8'hef;
      17'd25494: data = 8'hef;
      17'd25495: data = 8'hf1;
      17'd25496: data = 8'hf1;
      17'd25497: data = 8'hf2;
      17'd25498: data = 8'hf2;
      17'd25499: data = 8'hf4;
      17'd25500: data = 8'hf4;
      17'd25501: data = 8'hf4;
      17'd25502: data = 8'hf6;
      17'd25503: data = 8'hfa;
      17'd25504: data = 8'hfa;
      17'd25505: data = 8'hfa;
      17'd25506: data = 8'hf5;
      17'd25507: data = 8'hf4;
      17'd25508: data = 8'hf4;
      17'd25509: data = 8'hf2;
      17'd25510: data = 8'hed;
      17'd25511: data = 8'hef;
      17'd25512: data = 8'hef;
      17'd25513: data = 8'hf1;
      17'd25514: data = 8'hed;
      17'd25515: data = 8'he9;
      17'd25516: data = 8'he9;
      17'd25517: data = 8'hed;
      17'd25518: data = 8'hef;
      17'd25519: data = 8'hec;
      17'd25520: data = 8'hed;
      17'd25521: data = 8'hf2;
      17'd25522: data = 8'hf2;
      17'd25523: data = 8'hef;
      17'd25524: data = 8'hed;
      17'd25525: data = 8'hec;
      17'd25526: data = 8'he9;
      17'd25527: data = 8'he9;
      17'd25528: data = 8'hec;
      17'd25529: data = 8'heb;
      17'd25530: data = 8'he7;
      17'd25531: data = 8'he5;
      17'd25532: data = 8'he7;
      17'd25533: data = 8'he7;
      17'd25534: data = 8'he3;
      17'd25535: data = 8'he2;
      17'd25536: data = 8'he5;
      17'd25537: data = 8'he7;
      17'd25538: data = 8'he4;
      17'd25539: data = 8'he4;
      17'd25540: data = 8'he3;
      17'd25541: data = 8'he2;
      17'd25542: data = 8'he0;
      17'd25543: data = 8'he4;
      17'd25544: data = 8'he7;
      17'd25545: data = 8'he7;
      17'd25546: data = 8'heb;
      17'd25547: data = 8'hef;
      17'd25548: data = 8'hf4;
      17'd25549: data = 8'hf4;
      17'd25550: data = 8'hf1;
      17'd25551: data = 8'hf6;
      17'd25552: data = 8'hfc;
      17'd25553: data = 8'hfc;
      17'd25554: data = 8'hfd;
      17'd25555: data = 8'h00;
      17'd25556: data = 8'h01;
      17'd25557: data = 8'h02;
      17'd25558: data = 8'h01;
      17'd25559: data = 8'h02;
      17'd25560: data = 8'h05;
      17'd25561: data = 8'h09;
      17'd25562: data = 8'h0c;
      17'd25563: data = 8'h0d;
      17'd25564: data = 8'h0e;
      17'd25565: data = 8'h0e;
      17'd25566: data = 8'h0e;
      17'd25567: data = 8'h0e;
      17'd25568: data = 8'h0e;
      17'd25569: data = 8'h11;
      17'd25570: data = 8'h0e;
      17'd25571: data = 8'h12;
      17'd25572: data = 8'h15;
      17'd25573: data = 8'h16;
      17'd25574: data = 8'h15;
      17'd25575: data = 8'h15;
      17'd25576: data = 8'h16;
      17'd25577: data = 8'h16;
      17'd25578: data = 8'h15;
      17'd25579: data = 8'h15;
      17'd25580: data = 8'h16;
      17'd25581: data = 8'h15;
      17'd25582: data = 8'h13;
      17'd25583: data = 8'h13;
      17'd25584: data = 8'h0e;
      17'd25585: data = 8'h0d;
      17'd25586: data = 8'h0c;
      17'd25587: data = 8'h06;
      17'd25588: data = 8'h0a;
      17'd25589: data = 8'h0d;
      17'd25590: data = 8'h0c;
      17'd25591: data = 8'h0a;
      17'd25592: data = 8'h0d;
      17'd25593: data = 8'h0d;
      17'd25594: data = 8'h0c;
      17'd25595: data = 8'h0c;
      17'd25596: data = 8'h0c;
      17'd25597: data = 8'h0a;
      17'd25598: data = 8'h0c;
      17'd25599: data = 8'h0a;
      17'd25600: data = 8'h04;
      17'd25601: data = 8'h01;
      17'd25602: data = 8'h00;
      17'd25603: data = 8'hfe;
      17'd25604: data = 8'hfe;
      17'd25605: data = 8'hfe;
      17'd25606: data = 8'hfe;
      17'd25607: data = 8'hfe;
      17'd25608: data = 8'hfd;
      17'd25609: data = 8'hfe;
      17'd25610: data = 8'hfd;
      17'd25611: data = 8'hf9;
      17'd25612: data = 8'hfe;
      17'd25613: data = 8'h04;
      17'd25614: data = 8'h06;
      17'd25615: data = 8'h0c;
      17'd25616: data = 8'h0c;
      17'd25617: data = 8'h09;
      17'd25618: data = 8'h06;
      17'd25619: data = 8'h0c;
      17'd25620: data = 8'h0d;
      17'd25621: data = 8'h09;
      17'd25622: data = 8'h0e;
      17'd25623: data = 8'h13;
      17'd25624: data = 8'h13;
      17'd25625: data = 8'h11;
      17'd25626: data = 8'h0c;
      17'd25627: data = 8'h09;
      17'd25628: data = 8'h09;
      17'd25629: data = 8'h09;
      17'd25630: data = 8'h09;
      17'd25631: data = 8'h0c;
      17'd25632: data = 8'h0c;
      17'd25633: data = 8'h0a;
      17'd25634: data = 8'h0c;
      17'd25635: data = 8'h0a;
      17'd25636: data = 8'h06;
      17'd25637: data = 8'h05;
      17'd25638: data = 8'h09;
      17'd25639: data = 8'h0a;
      17'd25640: data = 8'h09;
      17'd25641: data = 8'h06;
      17'd25642: data = 8'h04;
      17'd25643: data = 8'h04;
      17'd25644: data = 8'h02;
      17'd25645: data = 8'hfd;
      17'd25646: data = 8'hfd;
      17'd25647: data = 8'hfd;
      17'd25648: data = 8'hfc;
      17'd25649: data = 8'hf9;
      17'd25650: data = 8'hf6;
      17'd25651: data = 8'hf2;
      17'd25652: data = 8'hef;
      17'd25653: data = 8'hef;
      17'd25654: data = 8'hec;
      17'd25655: data = 8'heb;
      17'd25656: data = 8'he9;
      17'd25657: data = 8'heb;
      17'd25658: data = 8'heb;
      17'd25659: data = 8'hec;
      17'd25660: data = 8'hec;
      17'd25661: data = 8'hed;
      17'd25662: data = 8'hf1;
      17'd25663: data = 8'hf1;
      17'd25664: data = 8'hef;
      17'd25665: data = 8'hf2;
      17'd25666: data = 8'hf6;
      17'd25667: data = 8'hfa;
      17'd25668: data = 8'hfc;
      17'd25669: data = 8'hfe;
      17'd25670: data = 8'hfe;
      17'd25671: data = 8'h00;
      17'd25672: data = 8'h01;
      17'd25673: data = 8'h01;
      17'd25674: data = 8'h02;
      17'd25675: data = 8'h02;
      17'd25676: data = 8'h02;
      17'd25677: data = 8'h04;
      17'd25678: data = 8'h06;
      17'd25679: data = 8'h06;
      17'd25680: data = 8'h05;
      17'd25681: data = 8'h09;
      17'd25682: data = 8'h09;
      17'd25683: data = 8'h0d;
      17'd25684: data = 8'h11;
      17'd25685: data = 8'h15;
      17'd25686: data = 8'h19;
      17'd25687: data = 8'h1a;
      17'd25688: data = 8'h1b;
      17'd25689: data = 8'h1b;
      17'd25690: data = 8'h24;
      17'd25691: data = 8'h1e;
      17'd25692: data = 8'h0a;
      17'd25693: data = 8'h13;
      17'd25694: data = 8'h1b;
      17'd25695: data = 8'h11;
      17'd25696: data = 8'h0e;
      17'd25697: data = 8'h15;
      17'd25698: data = 8'h11;
      17'd25699: data = 8'h06;
      17'd25700: data = 8'h06;
      17'd25701: data = 8'h0e;
      17'd25702: data = 8'h0c;
      17'd25703: data = 8'h05;
      17'd25704: data = 8'h0a;
      17'd25705: data = 8'h0e;
      17'd25706: data = 8'h09;
      17'd25707: data = 8'h05;
      17'd25708: data = 8'h05;
      17'd25709: data = 8'h02;
      17'd25710: data = 8'h05;
      17'd25711: data = 8'h06;
      17'd25712: data = 8'h04;
      17'd25713: data = 8'hfc;
      17'd25714: data = 8'h00;
      17'd25715: data = 8'h01;
      17'd25716: data = 8'hfa;
      17'd25717: data = 8'hfa;
      17'd25718: data = 8'hfc;
      17'd25719: data = 8'hf6;
      17'd25720: data = 8'hf6;
      17'd25721: data = 8'hf9;
      17'd25722: data = 8'hf5;
      17'd25723: data = 8'hec;
      17'd25724: data = 8'he9;
      17'd25725: data = 8'hed;
      17'd25726: data = 8'hef;
      17'd25727: data = 8'hef;
      17'd25728: data = 8'hef;
      17'd25729: data = 8'hf2;
      17'd25730: data = 8'hf5;
      17'd25731: data = 8'hfc;
      17'd25732: data = 8'hf5;
      17'd25733: data = 8'he9;
      17'd25734: data = 8'hed;
      17'd25735: data = 8'hf6;
      17'd25736: data = 8'hf9;
      17'd25737: data = 8'hf1;
      17'd25738: data = 8'hf1;
      17'd25739: data = 8'hf5;
      17'd25740: data = 8'hf5;
      17'd25741: data = 8'hec;
      17'd25742: data = 8'he9;
      17'd25743: data = 8'hec;
      17'd25744: data = 8'he9;
      17'd25745: data = 8'hec;
      17'd25746: data = 8'hf4;
      17'd25747: data = 8'hf5;
      17'd25748: data = 8'hef;
      17'd25749: data = 8'hed;
      17'd25750: data = 8'hf1;
      17'd25751: data = 8'hf1;
      17'd25752: data = 8'heb;
      17'd25753: data = 8'he5;
      17'd25754: data = 8'hef;
      17'd25755: data = 8'hf5;
      17'd25756: data = 8'hf2;
      17'd25757: data = 8'heb;
      17'd25758: data = 8'hed;
      17'd25759: data = 8'hf1;
      17'd25760: data = 8'hef;
      17'd25761: data = 8'heb;
      17'd25762: data = 8'he9;
      17'd25763: data = 8'hed;
      17'd25764: data = 8'hed;
      17'd25765: data = 8'he9;
      17'd25766: data = 8'he5;
      17'd25767: data = 8'he2;
      17'd25768: data = 8'he0;
      17'd25769: data = 8'hde;
      17'd25770: data = 8'he2;
      17'd25771: data = 8'he2;
      17'd25772: data = 8'he2;
      17'd25773: data = 8'he2;
      17'd25774: data = 8'he4;
      17'd25775: data = 8'he5;
      17'd25776: data = 8'he2;
      17'd25777: data = 8'he2;
      17'd25778: data = 8'he4;
      17'd25779: data = 8'heb;
      17'd25780: data = 8'heb;
      17'd25781: data = 8'hec;
      17'd25782: data = 8'hef;
      17'd25783: data = 8'hef;
      17'd25784: data = 8'hef;
      17'd25785: data = 8'hef;
      17'd25786: data = 8'hf1;
      17'd25787: data = 8'hf2;
      17'd25788: data = 8'hf4;
      17'd25789: data = 8'hf9;
      17'd25790: data = 8'hfa;
      17'd25791: data = 8'hfe;
      17'd25792: data = 8'h00;
      17'd25793: data = 8'h00;
      17'd25794: data = 8'h02;
      17'd25795: data = 8'h05;
      17'd25796: data = 8'h04;
      17'd25797: data = 8'h05;
      17'd25798: data = 8'h0c;
      17'd25799: data = 8'h0e;
      17'd25800: data = 8'h0d;
      17'd25801: data = 8'h0e;
      17'd25802: data = 8'h13;
      17'd25803: data = 8'h12;
      17'd25804: data = 8'h12;
      17'd25805: data = 8'h15;
      17'd25806: data = 8'h16;
      17'd25807: data = 8'h19;
      17'd25808: data = 8'h1a;
      17'd25809: data = 8'h19;
      17'd25810: data = 8'h16;
      17'd25811: data = 8'h16;
      17'd25812: data = 8'h1a;
      17'd25813: data = 8'h19;
      17'd25814: data = 8'h15;
      17'd25815: data = 8'h16;
      17'd25816: data = 8'h16;
      17'd25817: data = 8'h19;
      17'd25818: data = 8'h16;
      17'd25819: data = 8'h15;
      17'd25820: data = 8'h13;
      17'd25821: data = 8'h11;
      17'd25822: data = 8'h12;
      17'd25823: data = 8'h11;
      17'd25824: data = 8'h0a;
      17'd25825: data = 8'h0a;
      17'd25826: data = 8'h0e;
      17'd25827: data = 8'h0c;
      17'd25828: data = 8'h06;
      17'd25829: data = 8'h09;
      17'd25830: data = 8'h0c;
      17'd25831: data = 8'h0d;
      17'd25832: data = 8'h0c;
      17'd25833: data = 8'h0d;
      17'd25834: data = 8'h0d;
      17'd25835: data = 8'h09;
      17'd25836: data = 8'h02;
      17'd25837: data = 8'h01;
      17'd25838: data = 8'h01;
      17'd25839: data = 8'h01;
      17'd25840: data = 8'h00;
      17'd25841: data = 8'h01;
      17'd25842: data = 8'h00;
      17'd25843: data = 8'hfa;
      17'd25844: data = 8'hf5;
      17'd25845: data = 8'hf6;
      17'd25846: data = 8'hfd;
      17'd25847: data = 8'h00;
      17'd25848: data = 8'h02;
      17'd25849: data = 8'h0c;
      17'd25850: data = 8'h11;
      17'd25851: data = 8'h0d;
      17'd25852: data = 8'h0c;
      17'd25853: data = 8'h09;
      17'd25854: data = 8'h0e;
      17'd25855: data = 8'h11;
      17'd25856: data = 8'h0d;
      17'd25857: data = 8'h0e;
      17'd25858: data = 8'h15;
      17'd25859: data = 8'h11;
      17'd25860: data = 8'h06;
      17'd25861: data = 8'h05;
      17'd25862: data = 8'h05;
      17'd25863: data = 8'h04;
      17'd25864: data = 8'h04;
      17'd25865: data = 8'h09;
      17'd25866: data = 8'h0a;
      17'd25867: data = 8'h0a;
      17'd25868: data = 8'h0a;
      17'd25869: data = 8'h0d;
      17'd25870: data = 8'h0d;
      17'd25871: data = 8'h0a;
      17'd25872: data = 8'h09;
      17'd25873: data = 8'h0c;
      17'd25874: data = 8'h0d;
      17'd25875: data = 8'h0a;
      17'd25876: data = 8'h06;
      17'd25877: data = 8'h05;
      17'd25878: data = 8'h04;
      17'd25879: data = 8'h00;
      17'd25880: data = 8'hfd;
      17'd25881: data = 8'hfa;
      17'd25882: data = 8'hf9;
      17'd25883: data = 8'hf6;
      17'd25884: data = 8'hf5;
      17'd25885: data = 8'hf5;
      17'd25886: data = 8'hf5;
      17'd25887: data = 8'hf2;
      17'd25888: data = 8'hf2;
      17'd25889: data = 8'hf2;
      17'd25890: data = 8'hef;
      17'd25891: data = 8'hed;
      17'd25892: data = 8'hef;
      17'd25893: data = 8'hf2;
      17'd25894: data = 8'hf2;
      17'd25895: data = 8'hef;
      17'd25896: data = 8'hec;
      17'd25897: data = 8'hed;
      17'd25898: data = 8'hed;
      17'd25899: data = 8'hed;
      17'd25900: data = 8'hef;
      17'd25901: data = 8'hf5;
      17'd25902: data = 8'hfc;
      17'd25903: data = 8'hfd;
      17'd25904: data = 8'hfd;
      17'd25905: data = 8'hfd;
      17'd25906: data = 8'hfe;
      17'd25907: data = 8'hfe;
      17'd25908: data = 8'hfd;
      17'd25909: data = 8'hfe;
      17'd25910: data = 8'h01;
      17'd25911: data = 8'h02;
      17'd25912: data = 8'h04;
      17'd25913: data = 8'h05;
      17'd25914: data = 8'h06;
      17'd25915: data = 8'h06;
      17'd25916: data = 8'h06;
      17'd25917: data = 8'h0c;
      17'd25918: data = 8'h0e;
      17'd25919: data = 8'h0d;
      17'd25920: data = 8'h11;
      17'd25921: data = 8'h15;
      17'd25922: data = 8'h19;
      17'd25923: data = 8'h19;
      17'd25924: data = 8'h19;
      17'd25925: data = 8'h19;
      17'd25926: data = 8'h16;
      17'd25927: data = 8'h19;
      17'd25928: data = 8'h16;
      17'd25929: data = 8'h1a;
      17'd25930: data = 8'h1a;
      17'd25931: data = 8'h19;
      17'd25932: data = 8'h13;
      17'd25933: data = 8'h13;
      17'd25934: data = 8'h12;
      17'd25935: data = 8'h0d;
      17'd25936: data = 8'h0d;
      17'd25937: data = 8'h0e;
      17'd25938: data = 8'h0e;
      17'd25939: data = 8'h11;
      17'd25940: data = 8'h0e;
      17'd25941: data = 8'h11;
      17'd25942: data = 8'h0e;
      17'd25943: data = 8'h0d;
      17'd25944: data = 8'h0c;
      17'd25945: data = 8'h0a;
      17'd25946: data = 8'h06;
      17'd25947: data = 8'h04;
      17'd25948: data = 8'h02;
      17'd25949: data = 8'h00;
      17'd25950: data = 8'hfd;
      17'd25951: data = 8'hfc;
      17'd25952: data = 8'hfa;
      17'd25953: data = 8'hf9;
      17'd25954: data = 8'hf6;
      17'd25955: data = 8'hf5;
      17'd25956: data = 8'hf4;
      17'd25957: data = 8'hf4;
      17'd25958: data = 8'hf4;
      17'd25959: data = 8'hf4;
      17'd25960: data = 8'hf4;
      17'd25961: data = 8'hf4;
      17'd25962: data = 8'hf5;
      17'd25963: data = 8'hf6;
      17'd25964: data = 8'hf6;
      17'd25965: data = 8'hf6;
      17'd25966: data = 8'hf5;
      17'd25967: data = 8'hf2;
      17'd25968: data = 8'hf2;
      17'd25969: data = 8'hf1;
      17'd25970: data = 8'hed;
      17'd25971: data = 8'hef;
      17'd25972: data = 8'hed;
      17'd25973: data = 8'hec;
      17'd25974: data = 8'hed;
      17'd25975: data = 8'hed;
      17'd25976: data = 8'hed;
      17'd25977: data = 8'hf1;
      17'd25978: data = 8'hf2;
      17'd25979: data = 8'hef;
      17'd25980: data = 8'hed;
      17'd25981: data = 8'hed;
      17'd25982: data = 8'hed;
      17'd25983: data = 8'hed;
      17'd25984: data = 8'hed;
      17'd25985: data = 8'hed;
      17'd25986: data = 8'hef;
      17'd25987: data = 8'hf2;
      17'd25988: data = 8'hf2;
      17'd25989: data = 8'hf1;
      17'd25990: data = 8'hef;
      17'd25991: data = 8'hf1;
      17'd25992: data = 8'hef;
      17'd25993: data = 8'hec;
      17'd25994: data = 8'heb;
      17'd25995: data = 8'heb;
      17'd25996: data = 8'hec;
      17'd25997: data = 8'he9;
      17'd25998: data = 8'he9;
      17'd25999: data = 8'he5;
      17'd26000: data = 8'he5;
      17'd26001: data = 8'he5;
      17'd26002: data = 8'he5;
      17'd26003: data = 8'he5;
      17'd26004: data = 8'he4;
      17'd26005: data = 8'he4;
      17'd26006: data = 8'he3;
      17'd26007: data = 8'he4;
      17'd26008: data = 8'he2;
      17'd26009: data = 8'hdc;
      17'd26010: data = 8'he0;
      17'd26011: data = 8'he3;
      17'd26012: data = 8'he3;
      17'd26013: data = 8'he5;
      17'd26014: data = 8'he9;
      17'd26015: data = 8'hed;
      17'd26016: data = 8'hf1;
      17'd26017: data = 8'hef;
      17'd26018: data = 8'hef;
      17'd26019: data = 8'hf2;
      17'd26020: data = 8'hf2;
      17'd26021: data = 8'hf5;
      17'd26022: data = 8'hf5;
      17'd26023: data = 8'hf6;
      17'd26024: data = 8'hf9;
      17'd26025: data = 8'hfa;
      17'd26026: data = 8'hfa;
      17'd26027: data = 8'hfa;
      17'd26028: data = 8'hfd;
      17'd26029: data = 8'h00;
      17'd26030: data = 8'h01;
      17'd26031: data = 8'h01;
      17'd26032: data = 8'h04;
      17'd26033: data = 8'h05;
      17'd26034: data = 8'h06;
      17'd26035: data = 8'h0c;
      17'd26036: data = 8'h0c;
      17'd26037: data = 8'h0c;
      17'd26038: data = 8'h0d;
      17'd26039: data = 8'h12;
      17'd26040: data = 8'h13;
      17'd26041: data = 8'h13;
      17'd26042: data = 8'h15;
      17'd26043: data = 8'h16;
      17'd26044: data = 8'h19;
      17'd26045: data = 8'h16;
      17'd26046: data = 8'h15;
      17'd26047: data = 8'h16;
      17'd26048: data = 8'h19;
      17'd26049: data = 8'h19;
      17'd26050: data = 8'h16;
      17'd26051: data = 8'h15;
      17'd26052: data = 8'h15;
      17'd26053: data = 8'h13;
      17'd26054: data = 8'h15;
      17'd26055: data = 8'h15;
      17'd26056: data = 8'h15;
      17'd26057: data = 8'h15;
      17'd26058: data = 8'h13;
      17'd26059: data = 8'h16;
      17'd26060: data = 8'h15;
      17'd26061: data = 8'h13;
      17'd26062: data = 8'h12;
      17'd26063: data = 8'h12;
      17'd26064: data = 8'h0d;
      17'd26065: data = 8'h0d;
      17'd26066: data = 8'h11;
      17'd26067: data = 8'h0d;
      17'd26068: data = 8'h0c;
      17'd26069: data = 8'h0d;
      17'd26070: data = 8'h0e;
      17'd26071: data = 8'h0c;
      17'd26072: data = 8'h06;
      17'd26073: data = 8'h05;
      17'd26074: data = 8'h06;
      17'd26075: data = 8'h04;
      17'd26076: data = 8'h01;
      17'd26077: data = 8'h02;
      17'd26078: data = 8'h01;
      17'd26079: data = 8'hfd;
      17'd26080: data = 8'hfa;
      17'd26081: data = 8'hf9;
      17'd26082: data = 8'hf4;
      17'd26083: data = 8'hf2;
      17'd26084: data = 8'hf6;
      17'd26085: data = 8'hfe;
      17'd26086: data = 8'h02;
      17'd26087: data = 8'h01;
      17'd26088: data = 8'h02;
      17'd26089: data = 8'h05;
      17'd26090: data = 8'h09;
      17'd26091: data = 8'h06;
      17'd26092: data = 8'h05;
      17'd26093: data = 8'h06;
      17'd26094: data = 8'h09;
      17'd26095: data = 8'h0c;
      17'd26096: data = 8'h0a;
      17'd26097: data = 8'h05;
      17'd26098: data = 8'h02;
      17'd26099: data = 8'h01;
      17'd26100: data = 8'h02;
      17'd26101: data = 8'h04;
      17'd26102: data = 8'h02;
      17'd26103: data = 8'h04;
      17'd26104: data = 8'h09;
      17'd26105: data = 8'h0c;
      17'd26106: data = 8'h0d;
      17'd26107: data = 8'h0c;
      17'd26108: data = 8'h0a;
      17'd26109: data = 8'h09;
      17'd26110: data = 8'h0a;
      17'd26111: data = 8'h0a;
      17'd26112: data = 8'h06;
      17'd26113: data = 8'h04;
      17'd26114: data = 8'h05;
      17'd26115: data = 8'h06;
      17'd26116: data = 8'h04;
      17'd26117: data = 8'h00;
      17'd26118: data = 8'h01;
      17'd26119: data = 8'h01;
      17'd26120: data = 8'h00;
      17'd26121: data = 8'hfe;
      17'd26122: data = 8'hfd;
      17'd26123: data = 8'hfc;
      17'd26124: data = 8'hf9;
      17'd26125: data = 8'hf5;
      17'd26126: data = 8'hf4;
      17'd26127: data = 8'hf1;
      17'd26128: data = 8'hef;
      17'd26129: data = 8'hef;
      17'd26130: data = 8'hf1;
      17'd26131: data = 8'hef;
      17'd26132: data = 8'hef;
      17'd26133: data = 8'hf1;
      17'd26134: data = 8'hf1;
      17'd26135: data = 8'hf1;
      17'd26136: data = 8'hef;
      17'd26137: data = 8'hf1;
      17'd26138: data = 8'hf2;
      17'd26139: data = 8'hf2;
      17'd26140: data = 8'hf5;
      17'd26141: data = 8'hf5;
      17'd26142: data = 8'hf5;
      17'd26143: data = 8'hf9;
      17'd26144: data = 8'hfa;
      17'd26145: data = 8'hfa;
      17'd26146: data = 8'hfc;
      17'd26147: data = 8'hfc;
      17'd26148: data = 8'hfc;
      17'd26149: data = 8'hfe;
      17'd26150: data = 8'h00;
      17'd26151: data = 8'h01;
      17'd26152: data = 8'h01;
      17'd26153: data = 8'h02;
      17'd26154: data = 8'h04;
      17'd26155: data = 8'h06;
      17'd26156: data = 8'h09;
      17'd26157: data = 8'h0c;
      17'd26158: data = 8'h11;
      17'd26159: data = 8'h11;
      17'd26160: data = 8'h12;
      17'd26161: data = 8'h15;
      17'd26162: data = 8'h15;
      17'd26163: data = 8'h15;
      17'd26164: data = 8'h13;
      17'd26165: data = 8'h12;
      17'd26166: data = 8'h12;
      17'd26167: data = 8'h13;
      17'd26168: data = 8'h12;
      17'd26169: data = 8'h11;
      17'd26170: data = 8'h12;
      17'd26171: data = 8'h13;
      17'd26172: data = 8'h13;
      17'd26173: data = 8'h13;
      17'd26174: data = 8'h13;
      17'd26175: data = 8'h11;
      17'd26176: data = 8'h0e;
      17'd26177: data = 8'h0d;
      17'd26178: data = 8'h0d;
      17'd26179: data = 8'h0a;
      17'd26180: data = 8'h06;
      17'd26181: data = 8'h06;
      17'd26182: data = 8'h05;
      17'd26183: data = 8'h02;
      17'd26184: data = 8'h01;
      17'd26185: data = 8'h00;
      17'd26186: data = 8'hfe;
      17'd26187: data = 8'hfe;
      17'd26188: data = 8'hfd;
      17'd26189: data = 8'hfd;
      17'd26190: data = 8'hfc;
      17'd26191: data = 8'hfc;
      17'd26192: data = 8'hfc;
      17'd26193: data = 8'hf9;
      17'd26194: data = 8'hf6;
      17'd26195: data = 8'hf6;
      17'd26196: data = 8'hf6;
      17'd26197: data = 8'hf5;
      17'd26198: data = 8'hf2;
      17'd26199: data = 8'hf1;
      17'd26200: data = 8'hef;
      17'd26201: data = 8'hef;
      17'd26202: data = 8'hed;
      17'd26203: data = 8'hed;
      17'd26204: data = 8'hf1;
      17'd26205: data = 8'hf4;
      17'd26206: data = 8'hf4;
      17'd26207: data = 8'hfa;
      17'd26208: data = 8'he7;
      17'd26209: data = 8'he9;
      17'd26210: data = 8'hfd;
      17'd26211: data = 8'hf5;
      17'd26212: data = 8'hed;
      17'd26213: data = 8'hf2;
      17'd26214: data = 8'hfa;
      17'd26215: data = 8'hf2;
      17'd26216: data = 8'he9;
      17'd26217: data = 8'hf5;
      17'd26218: data = 8'hf2;
      17'd26219: data = 8'he3;
      17'd26220: data = 8'hec;
      17'd26221: data = 8'hf6;
      17'd26222: data = 8'hf1;
      17'd26223: data = 8'hec;
      17'd26224: data = 8'hef;
      17'd26225: data = 8'he9;
      17'd26226: data = 8'heb;
      17'd26227: data = 8'hec;
      17'd26228: data = 8'he3;
      17'd26229: data = 8'he2;
      17'd26230: data = 8'hed;
      17'd26231: data = 8'hed;
      17'd26232: data = 8'he5;
      17'd26233: data = 8'hef;
      17'd26234: data = 8'hf6;
      17'd26235: data = 8'hed;
      17'd26236: data = 8'he7;
      17'd26237: data = 8'hef;
      17'd26238: data = 8'heb;
      17'd26239: data = 8'he3;
      17'd26240: data = 8'he7;
      17'd26241: data = 8'heb;
      17'd26242: data = 8'he4;
      17'd26243: data = 8'he7;
      17'd26244: data = 8'hec;
      17'd26245: data = 8'he9;
      17'd26246: data = 8'he7;
      17'd26247: data = 8'hec;
      17'd26248: data = 8'hed;
      17'd26249: data = 8'hef;
      17'd26250: data = 8'hf2;
      17'd26251: data = 8'hf2;
      17'd26252: data = 8'hf2;
      17'd26253: data = 8'hf1;
      17'd26254: data = 8'hef;
      17'd26255: data = 8'hf1;
      17'd26256: data = 8'hf2;
      17'd26257: data = 8'hf4;
      17'd26258: data = 8'hf4;
      17'd26259: data = 8'hfa;
      17'd26260: data = 8'hfe;
      17'd26261: data = 8'hfc;
      17'd26262: data = 8'hfc;
      17'd26263: data = 8'h01;
      17'd26264: data = 8'h01;
      17'd26265: data = 8'h01;
      17'd26266: data = 8'hf4;
      17'd26267: data = 8'he9;
      17'd26268: data = 8'hed;
      17'd26269: data = 8'hfa;
      17'd26270: data = 8'h04;
      17'd26271: data = 8'h02;
      17'd26272: data = 8'h00;
      17'd26273: data = 8'h06;
      17'd26274: data = 8'h09;
      17'd26275: data = 8'h11;
      17'd26276: data = 8'h19;
      17'd26277: data = 8'h15;
      17'd26278: data = 8'h15;
      17'd26279: data = 8'h1a;
      17'd26280: data = 8'h1c;
      17'd26281: data = 8'h19;
      17'd26282: data = 8'h0e;
      17'd26283: data = 8'h0a;
      17'd26284: data = 8'h12;
      17'd26285: data = 8'h16;
      17'd26286: data = 8'h19;
      17'd26287: data = 8'h0d;
      17'd26288: data = 8'h0c;
      17'd26289: data = 8'h12;
      17'd26290: data = 8'h16;
      17'd26291: data = 8'h15;
      17'd26292: data = 8'h16;
      17'd26293: data = 8'h19;
      17'd26294: data = 8'h15;
      17'd26295: data = 8'h11;
      17'd26296: data = 8'h15;
      17'd26297: data = 8'h19;
      17'd26298: data = 8'h12;
      17'd26299: data = 8'h16;
      17'd26300: data = 8'h16;
      17'd26301: data = 8'h0e;
      17'd26302: data = 8'h0a;
      17'd26303: data = 8'h11;
      17'd26304: data = 8'h15;
      17'd26305: data = 8'h15;
      17'd26306: data = 8'h0e;
      17'd26307: data = 8'h13;
      17'd26308: data = 8'h13;
      17'd26309: data = 8'h06;
      17'd26310: data = 8'hf6;
      17'd26311: data = 8'hf1;
      17'd26312: data = 8'hf2;
      17'd26313: data = 8'hf5;
      17'd26314: data = 8'hfd;
      17'd26315: data = 8'h04;
      17'd26316: data = 8'h05;
      17'd26317: data = 8'h02;
      17'd26318: data = 8'h05;
      17'd26319: data = 8'h00;
      17'd26320: data = 8'hf9;
      17'd26321: data = 8'hfa;
      17'd26322: data = 8'h09;
      17'd26323: data = 8'h13;
      17'd26324: data = 8'h0e;
      17'd26325: data = 8'h0a;
      17'd26326: data = 8'h0d;
      17'd26327: data = 8'h11;
      17'd26328: data = 8'h0c;
      17'd26329: data = 8'h01;
      17'd26330: data = 8'h02;
      17'd26331: data = 8'h05;
      17'd26332: data = 8'h0c;
      17'd26333: data = 8'h1a;
      17'd26334: data = 8'h1c;
      17'd26335: data = 8'h15;
      17'd26336: data = 8'h16;
      17'd26337: data = 8'h1c;
      17'd26338: data = 8'h15;
      17'd26339: data = 8'h05;
      17'd26340: data = 8'hfe;
      17'd26341: data = 8'h05;
      17'd26342: data = 8'h11;
      17'd26343: data = 8'h11;
      17'd26344: data = 8'h0a;
      17'd26345: data = 8'h09;
      17'd26346: data = 8'h05;
      17'd26347: data = 8'h01;
      17'd26348: data = 8'hfc;
      17'd26349: data = 8'hfd;
      17'd26350: data = 8'h00;
      17'd26351: data = 8'h06;
      17'd26352: data = 8'h11;
      17'd26353: data = 8'h0d;
      17'd26354: data = 8'h01;
      17'd26355: data = 8'hfe;
      17'd26356: data = 8'hfc;
      17'd26357: data = 8'hf1;
      17'd26358: data = 8'he7;
      17'd26359: data = 8'he5;
      17'd26360: data = 8'he5;
      17'd26361: data = 8'he5;
      17'd26362: data = 8'he3;
      17'd26363: data = 8'he0;
      17'd26364: data = 8'he3;
      17'd26365: data = 8'he2;
      17'd26366: data = 8'he3;
      17'd26367: data = 8'he5;
      17'd26368: data = 8'he7;
      17'd26369: data = 8'heb;
      17'd26370: data = 8'hf5;
      17'd26371: data = 8'hfe;
      17'd26372: data = 8'hfd;
      17'd26373: data = 8'hf6;
      17'd26374: data = 8'hfa;
      17'd26375: data = 8'hf9;
      17'd26376: data = 8'hed;
      17'd26377: data = 8'he9;
      17'd26378: data = 8'hf1;
      17'd26379: data = 8'hfc;
      17'd26380: data = 8'h00;
      17'd26381: data = 8'h05;
      17'd26382: data = 8'h06;
      17'd26383: data = 8'h05;
      17'd26384: data = 8'h09;
      17'd26385: data = 8'h0c;
      17'd26386: data = 8'h0d;
      17'd26387: data = 8'h12;
      17'd26388: data = 8'h1a;
      17'd26389: data = 8'h1c;
      17'd26390: data = 8'h1e;
      17'd26391: data = 8'h1a;
      17'd26392: data = 8'h15;
      17'd26393: data = 8'h13;
      17'd26394: data = 8'h11;
      17'd26395: data = 8'h0d;
      17'd26396: data = 8'h0e;
      17'd26397: data = 8'h12;
      17'd26398: data = 8'h16;
      17'd26399: data = 8'h1c;
      17'd26400: data = 8'h1e;
      17'd26401: data = 8'h23;
      17'd26402: data = 8'h26;
      17'd26403: data = 8'h1f;
      17'd26404: data = 8'h1b;
      17'd26405: data = 8'h16;
      17'd26406: data = 8'h13;
      17'd26407: data = 8'h16;
      17'd26408: data = 8'h19;
      17'd26409: data = 8'h12;
      17'd26410: data = 8'h0c;
      17'd26411: data = 8'h05;
      17'd26412: data = 8'hfd;
      17'd26413: data = 8'hf6;
      17'd26414: data = 8'hf5;
      17'd26415: data = 8'hfa;
      17'd26416: data = 8'h00;
      17'd26417: data = 8'h05;
      17'd26418: data = 8'h06;
      17'd26419: data = 8'h05;
      17'd26420: data = 8'h04;
      17'd26421: data = 8'h00;
      17'd26422: data = 8'hfd;
      17'd26423: data = 8'hf9;
      17'd26424: data = 8'hf6;
      17'd26425: data = 8'hf5;
      17'd26426: data = 8'hf9;
      17'd26427: data = 8'hf9;
      17'd26428: data = 8'hf5;
      17'd26429: data = 8'hf4;
      17'd26430: data = 8'hf2;
      17'd26431: data = 8'hf1;
      17'd26432: data = 8'hed;
      17'd26433: data = 8'hed;
      17'd26434: data = 8'hf1;
      17'd26435: data = 8'hfa;
      17'd26436: data = 8'h00;
      17'd26437: data = 8'h02;
      17'd26438: data = 8'h04;
      17'd26439: data = 8'h01;
      17'd26440: data = 8'hfa;
      17'd26441: data = 8'hf4;
      17'd26442: data = 8'hef;
      17'd26443: data = 8'hed;
      17'd26444: data = 8'hf4;
      17'd26445: data = 8'hf5;
      17'd26446: data = 8'hf4;
      17'd26447: data = 8'hf2;
      17'd26448: data = 8'hf5;
      17'd26449: data = 8'hf4;
      17'd26450: data = 8'hf5;
      17'd26451: data = 8'hf5;
      17'd26452: data = 8'hf5;
      17'd26453: data = 8'hf6;
      17'd26454: data = 8'hf6;
      17'd26455: data = 8'hf4;
      17'd26456: data = 8'hf1;
      17'd26457: data = 8'hed;
      17'd26458: data = 8'he9;
      17'd26459: data = 8'he3;
      17'd26460: data = 8'hdc;
      17'd26461: data = 8'hd6;
      17'd26462: data = 8'hd8;
      17'd26463: data = 8'he2;
      17'd26464: data = 8'he5;
      17'd26465: data = 8'he9;
      17'd26466: data = 8'heb;
      17'd26467: data = 8'he9;
      17'd26468: data = 8'he9;
      17'd26469: data = 8'heb;
      17'd26470: data = 8'he4;
      17'd26471: data = 8'he2;
      17'd26472: data = 8'he3;
      17'd26473: data = 8'he3;
      17'd26474: data = 8'he0;
      17'd26475: data = 8'hdc;
      17'd26476: data = 8'hda;
      17'd26477: data = 8'hdc;
      17'd26478: data = 8'he3;
      17'd26479: data = 8'he3;
      17'd26480: data = 8'he7;
      17'd26481: data = 8'hf1;
      17'd26482: data = 8'hf9;
      17'd26483: data = 8'hfd;
      17'd26484: data = 8'hfe;
      17'd26485: data = 8'hfe;
      17'd26486: data = 8'hfa;
      17'd26487: data = 8'hf5;
      17'd26488: data = 8'hf2;
      17'd26489: data = 8'hf2;
      17'd26490: data = 8'hf2;
      17'd26491: data = 8'hf5;
      17'd26492: data = 8'hfc;
      17'd26493: data = 8'h00;
      17'd26494: data = 8'h00;
      17'd26495: data = 8'h04;
      17'd26496: data = 8'h0c;
      17'd26497: data = 8'h0d;
      17'd26498: data = 8'h0e;
      17'd26499: data = 8'h11;
      17'd26500: data = 8'h16;
      17'd26501: data = 8'h16;
      17'd26502: data = 8'h12;
      17'd26503: data = 8'h0c;
      17'd26504: data = 8'h09;
      17'd26505: data = 8'h05;
      17'd26506: data = 8'h01;
      17'd26507: data = 8'h00;
      17'd26508: data = 8'h00;
      17'd26509: data = 8'h01;
      17'd26510: data = 8'h05;
      17'd26511: data = 8'h0e;
      17'd26512: data = 8'h12;
      17'd26513: data = 8'h12;
      17'd26514: data = 8'h11;
      17'd26515: data = 8'h12;
      17'd26516: data = 8'h12;
      17'd26517: data = 8'h0e;
      17'd26518: data = 8'h0c;
      17'd26519: data = 8'h0c;
      17'd26520: data = 8'h0e;
      17'd26521: data = 8'h0a;
      17'd26522: data = 8'h06;
      17'd26523: data = 8'h04;
      17'd26524: data = 8'h09;
      17'd26525: data = 8'h01;
      17'd26526: data = 8'h04;
      17'd26527: data = 8'h00;
      17'd26528: data = 8'h06;
      17'd26529: data = 8'h0a;
      17'd26530: data = 8'h0c;
      17'd26531: data = 8'h12;
      17'd26532: data = 8'h05;
      17'd26533: data = 8'h09;
      17'd26534: data = 8'h06;
      17'd26535: data = 8'h0c;
      17'd26536: data = 8'h01;
      17'd26537: data = 8'h09;
      17'd26538: data = 8'hfe;
      17'd26539: data = 8'h09;
      17'd26540: data = 8'h12;
      17'd26541: data = 8'h09;
      17'd26542: data = 8'h0a;
      17'd26543: data = 8'h12;
      17'd26544: data = 8'h0c;
      17'd26545: data = 8'hf6;
      17'd26546: data = 8'hfe;
      17'd26547: data = 8'heb;
      17'd26548: data = 8'he4;
      17'd26549: data = 8'he3;
      17'd26550: data = 8'hef;
      17'd26551: data = 8'hec;
      17'd26552: data = 8'he4;
      17'd26553: data = 8'he5;
      17'd26554: data = 8'hf6;
      17'd26555: data = 8'hf9;
      17'd26556: data = 8'hfd;
      17'd26557: data = 8'h12;
      17'd26558: data = 8'h23;
      17'd26559: data = 8'h22;
      17'd26560: data = 8'h13;
      17'd26561: data = 8'h1b;
      17'd26562: data = 8'h11;
      17'd26563: data = 8'h04;
      17'd26564: data = 8'hfc;
      17'd26565: data = 8'h0e;
      17'd26566: data = 8'h0e;
      17'd26567: data = 8'h09;
      17'd26568: data = 8'h0c;
      17'd26569: data = 8'h19;
      17'd26570: data = 8'h1c;
      17'd26571: data = 8'h1f;
      17'd26572: data = 8'h27;
      17'd26573: data = 8'h31;
      17'd26574: data = 8'h2b;
      17'd26575: data = 8'h1a;
      17'd26576: data = 8'h1e;
      17'd26577: data = 8'h1e;
      17'd26578: data = 8'h13;
      17'd26579: data = 8'h02;
      17'd26580: data = 8'h02;
      17'd26581: data = 8'hfa;
      17'd26582: data = 8'he7;
      17'd26583: data = 8'he3;
      17'd26584: data = 8'hf1;
      17'd26585: data = 8'hf6;
      17'd26586: data = 8'hfc;
      17'd26587: data = 8'h05;
      17'd26588: data = 8'h0d;
      17'd26589: data = 8'h04;
      17'd26590: data = 8'hfa;
      17'd26591: data = 8'hef;
      17'd26592: data = 8'hed;
      17'd26593: data = 8'he4;
      17'd26594: data = 8'he0;
      17'd26595: data = 8'hde;
      17'd26596: data = 8'hd6;
      17'd26597: data = 8'hcb;
      17'd26598: data = 8'hc6;
      17'd26599: data = 8'hd1;
      17'd26600: data = 8'hd2;
      17'd26601: data = 8'hdc;
      17'd26602: data = 8'heb;
      17'd26603: data = 8'hf2;
      17'd26604: data = 8'hf9;
      17'd26605: data = 8'hfd;
      17'd26606: data = 8'h00;
      17'd26607: data = 8'h06;
      17'd26608: data = 8'h04;
      17'd26609: data = 8'h01;
      17'd26610: data = 8'h02;
      17'd26611: data = 8'hfd;
      17'd26612: data = 8'hfd;
      17'd26613: data = 8'h05;
      17'd26614: data = 8'h0e;
      17'd26615: data = 8'h15;
      17'd26616: data = 8'h1c;
      17'd26617: data = 8'h24;
      17'd26618: data = 8'h27;
      17'd26619: data = 8'h26;
      17'd26620: data = 8'h26;
      17'd26621: data = 8'h2f;
      17'd26622: data = 8'h34;
      17'd26623: data = 8'h2f;
      17'd26624: data = 8'h2d;
      17'd26625: data = 8'h24;
      17'd26626: data = 8'h19;
      17'd26627: data = 8'h11;
      17'd26628: data = 8'h0e;
      17'd26629: data = 8'h12;
      17'd26630: data = 8'h16;
      17'd26631: data = 8'h1a;
      17'd26632: data = 8'h1f;
      17'd26633: data = 8'h1f;
      17'd26634: data = 8'h1a;
      17'd26635: data = 8'h19;
      17'd26636: data = 8'h1b;
      17'd26637: data = 8'h12;
      17'd26638: data = 8'h06;
      17'd26639: data = 8'hfe;
      17'd26640: data = 8'hf4;
      17'd26641: data = 8'hf1;
      17'd26642: data = 8'he7;
      17'd26643: data = 8'he4;
      17'd26644: data = 8'he5;
      17'd26645: data = 8'he5;
      17'd26646: data = 8'he3;
      17'd26647: data = 8'he4;
      17'd26648: data = 8'he5;
      17'd26649: data = 8'he7;
      17'd26650: data = 8'hf1;
      17'd26651: data = 8'hf6;
      17'd26652: data = 8'hf9;
      17'd26653: data = 8'hf2;
      17'd26654: data = 8'heb;
      17'd26655: data = 8'he4;
      17'd26656: data = 8'he3;
      17'd26657: data = 8'he2;
      17'd26658: data = 8'he9;
      17'd26659: data = 8'hf1;
      17'd26660: data = 8'hf5;
      17'd26661: data = 8'hfa;
      17'd26662: data = 8'h00;
      17'd26663: data = 8'h05;
      17'd26664: data = 8'h0a;
      17'd26665: data = 8'h13;
      17'd26666: data = 8'h16;
      17'd26667: data = 8'h16;
      17'd26668: data = 8'h15;
      17'd26669: data = 8'h11;
      17'd26670: data = 8'h0d;
      17'd26671: data = 8'h06;
      17'd26672: data = 8'h01;
      17'd26673: data = 8'h00;
      17'd26674: data = 8'hfd;
      17'd26675: data = 8'hf9;
      17'd26676: data = 8'hfd;
      17'd26677: data = 8'h01;
      17'd26678: data = 8'h05;
      17'd26679: data = 8'h0a;
      17'd26680: data = 8'h0a;
      17'd26681: data = 8'h06;
      17'd26682: data = 8'h02;
      17'd26683: data = 8'hf5;
      17'd26684: data = 8'heb;
      17'd26685: data = 8'he7;
      17'd26686: data = 8'he3;
      17'd26687: data = 8'he0;
      17'd26688: data = 8'he3;
      17'd26689: data = 8'hde;
      17'd26690: data = 8'hd5;
      17'd26691: data = 8'hd6;
      17'd26692: data = 8'hd6;
      17'd26693: data = 8'hd8;
      17'd26694: data = 8'hda;
      17'd26695: data = 8'hdc;
      17'd26696: data = 8'hdc;
      17'd26697: data = 8'hdc;
      17'd26698: data = 8'hd8;
      17'd26699: data = 8'hdb;
      17'd26700: data = 8'hda;
      17'd26701: data = 8'hd1;
      17'd26702: data = 8'hca;
      17'd26703: data = 8'hcd;
      17'd26704: data = 8'hd3;
      17'd26705: data = 8'hd8;
      17'd26706: data = 8'he3;
      17'd26707: data = 8'hed;
      17'd26708: data = 8'hf4;
      17'd26709: data = 8'hf6;
      17'd26710: data = 8'hf9;
      17'd26711: data = 8'hfa;
      17'd26712: data = 8'hf9;
      17'd26713: data = 8'hf9;
      17'd26714: data = 8'hfd;
      17'd26715: data = 8'hfe;
      17'd26716: data = 8'hfe;
      17'd26717: data = 8'hfa;
      17'd26718: data = 8'hfc;
      17'd26719: data = 8'h01;
      17'd26720: data = 8'h01;
      17'd26721: data = 8'h05;
      17'd26722: data = 8'h0d;
      17'd26723: data = 8'h11;
      17'd26724: data = 8'h11;
      17'd26725: data = 8'h12;
      17'd26726: data = 8'h12;
      17'd26727: data = 8'h0a;
      17'd26728: data = 8'h06;
      17'd26729: data = 8'h02;
      17'd26730: data = 8'hfd;
      17'd26731: data = 8'hfa;
      17'd26732: data = 8'hfa;
      17'd26733: data = 8'hfe;
      17'd26734: data = 8'h00;
      17'd26735: data = 8'h02;
      17'd26736: data = 8'h04;
      17'd26737: data = 8'h05;
      17'd26738: data = 8'h02;
      17'd26739: data = 8'h01;
      17'd26740: data = 8'h01;
      17'd26741: data = 8'hfe;
      17'd26742: data = 8'h01;
      17'd26743: data = 8'h00;
      17'd26744: data = 8'hfd;
      17'd26745: data = 8'hfa;
      17'd26746: data = 8'hf5;
      17'd26747: data = 8'hed;
      17'd26748: data = 8'heb;
      17'd26749: data = 8'hed;
      17'd26750: data = 8'hf1;
      17'd26751: data = 8'hf9;
      17'd26752: data = 8'hfc;
      17'd26753: data = 8'h02;
      17'd26754: data = 8'h04;
      17'd26755: data = 8'h05;
      17'd26756: data = 8'h04;
      17'd26757: data = 8'h04;
      17'd26758: data = 8'hfe;
      17'd26759: data = 8'hfd;
      17'd26760: data = 8'h05;
      17'd26761: data = 8'h02;
      17'd26762: data = 8'hfe;
      17'd26763: data = 8'h09;
      17'd26764: data = 8'h12;
      17'd26765: data = 8'h0e;
      17'd26766: data = 8'h1e;
      17'd26767: data = 8'h13;
      17'd26768: data = 8'h0a;
      17'd26769: data = 8'h15;
      17'd26770: data = 8'h19;
      17'd26771: data = 8'h16;
      17'd26772: data = 8'h1c;
      17'd26773: data = 8'h19;
      17'd26774: data = 8'h13;
      17'd26775: data = 8'h1f;
      17'd26776: data = 8'h13;
      17'd26777: data = 8'h0d;
      17'd26778: data = 8'h12;
      17'd26779: data = 8'h0e;
      17'd26780: data = 8'h11;
      17'd26781: data = 8'h0e;
      17'd26782: data = 8'hfd;
      17'd26783: data = 8'hfd;
      17'd26784: data = 8'h00;
      17'd26785: data = 8'heb;
      17'd26786: data = 8'hfc;
      17'd26787: data = 8'hf9;
      17'd26788: data = 8'he4;
      17'd26789: data = 8'he7;
      17'd26790: data = 8'hed;
      17'd26791: data = 8'he2;
      17'd26792: data = 8'hd5;
      17'd26793: data = 8'hca;
      17'd26794: data = 8'hde;
      17'd26795: data = 8'hfa;
      17'd26796: data = 8'hfa;
      17'd26797: data = 8'h19;
      17'd26798: data = 8'h34;
      17'd26799: data = 8'h26;
      17'd26800: data = 8'h1f;
      17'd26801: data = 8'h27;
      17'd26802: data = 8'h16;
      17'd26803: data = 8'h0e;
      17'd26804: data = 8'h0e;
      17'd26805: data = 8'h15;
      17'd26806: data = 8'h26;
      17'd26807: data = 8'h16;
      17'd26808: data = 8'h12;
      17'd26809: data = 8'h2b;
      17'd26810: data = 8'h2c;
      17'd26811: data = 8'h26;
      17'd26812: data = 8'h36;
      17'd26813: data = 8'h3e;
      17'd26814: data = 8'h3a;
      17'd26815: data = 8'h36;
      17'd26816: data = 8'h2d;
      17'd26817: data = 8'h2b;
      17'd26818: data = 8'h13;
      17'd26819: data = 8'hfa;
      17'd26820: data = 8'hf9;
      17'd26821: data = 8'he9;
      17'd26822: data = 8'hd1;
      17'd26823: data = 8'hda;
      17'd26824: data = 8'he7;
      17'd26825: data = 8'he9;
      17'd26826: data = 8'hed;
      17'd26827: data = 8'hf4;
      17'd26828: data = 8'hf5;
      17'd26829: data = 8'heb;
      17'd26830: data = 8'hd3;
      17'd26831: data = 8'hd6;
      17'd26832: data = 8'hd6;
      17'd26833: data = 8'hca;
      17'd26834: data = 8'hcd;
      17'd26835: data = 8'hcb;
      17'd26836: data = 8'hc0;
      17'd26837: data = 8'hbb;
      17'd26838: data = 8'hbb;
      17'd26839: data = 8'hc4;
      17'd26840: data = 8'hd1;
      17'd26841: data = 8'hdc;
      17'd26842: data = 8'hf2;
      17'd26843: data = 8'h02;
      17'd26844: data = 8'h02;
      17'd26845: data = 8'h05;
      17'd26846: data = 8'h0a;
      17'd26847: data = 8'h09;
      17'd26848: data = 8'h0d;
      17'd26849: data = 8'h09;
      17'd26850: data = 8'h0c;
      17'd26851: data = 8'h15;
      17'd26852: data = 8'h15;
      17'd26853: data = 8'h1f;
      17'd26854: data = 8'h31;
      17'd26855: data = 8'h33;
      17'd26856: data = 8'h3d;
      17'd26857: data = 8'h43;
      17'd26858: data = 8'h3d;
      17'd26859: data = 8'h3e;
      17'd26860: data = 8'h40;
      17'd26861: data = 8'h3d;
      17'd26862: data = 8'h42;
      17'd26863: data = 8'h35;
      17'd26864: data = 8'h26;
      17'd26865: data = 8'h1f;
      17'd26866: data = 8'h05;
      17'd26867: data = 8'h04;
      17'd26868: data = 8'h11;
      17'd26869: data = 8'h11;
      17'd26870: data = 8'h16;
      17'd26871: data = 8'h1b;
      17'd26872: data = 8'h15;
      17'd26873: data = 8'h0e;
      17'd26874: data = 8'h04;
      17'd26875: data = 8'hfc;
      17'd26876: data = 8'hfa;
      17'd26877: data = 8'he9;
      17'd26878: data = 8'he0;
      17'd26879: data = 8'hde;
      17'd26880: data = 8'hd1;
      17'd26881: data = 8'hcb;
      17'd26882: data = 8'hd2;
      17'd26883: data = 8'hd2;
      17'd26884: data = 8'hd8;
      17'd26885: data = 8'hdb;
      17'd26886: data = 8'hdc;
      17'd26887: data = 8'he5;
      17'd26888: data = 8'he9;
      17'd26889: data = 8'heb;
      17'd26890: data = 8'hf9;
      17'd26891: data = 8'hf5;
      17'd26892: data = 8'hef;
      17'd26893: data = 8'hf1;
      17'd26894: data = 8'he4;
      17'd26895: data = 8'he4;
      17'd26896: data = 8'hf1;
      17'd26897: data = 8'hf6;
      17'd26898: data = 8'h05;
      17'd26899: data = 8'h13;
      17'd26900: data = 8'h16;
      17'd26901: data = 8'h1f;
      17'd26902: data = 8'h1e;
      17'd26903: data = 8'h1a;
      17'd26904: data = 8'h1f;
      17'd26905: data = 8'h1f;
      17'd26906: data = 8'h1a;
      17'd26907: data = 8'h19;
      17'd26908: data = 8'h11;
      17'd26909: data = 8'h06;
      17'd26910: data = 8'h05;
      17'd26911: data = 8'hfe;
      17'd26912: data = 8'hfe;
      17'd26913: data = 8'h02;
      17'd26914: data = 8'hfe;
      17'd26915: data = 8'hfd;
      17'd26916: data = 8'hfd;
      17'd26917: data = 8'hfa;
      17'd26918: data = 8'hfe;
      17'd26919: data = 8'hfc;
      17'd26920: data = 8'hef;
      17'd26921: data = 8'he7;
      17'd26922: data = 8'hd3;
      17'd26923: data = 8'hc2;
      17'd26924: data = 8'hc6;
      17'd26925: data = 8'hc4;
      17'd26926: data = 8'hc5;
      17'd26927: data = 8'hd6;
      17'd26928: data = 8'hd5;
      17'd26929: data = 8'hd5;
      17'd26930: data = 8'hdb;
      17'd26931: data = 8'hd5;
      17'd26932: data = 8'hda;
      17'd26933: data = 8'he0;
      17'd26934: data = 8'hde;
      17'd26935: data = 8'heb;
      17'd26936: data = 8'he5;
      17'd26937: data = 8'hd8;
      17'd26938: data = 8'hde;
      17'd26939: data = 8'hde;
      17'd26940: data = 8'hdb;
      17'd26941: data = 8'he7;
      17'd26942: data = 8'hef;
      17'd26943: data = 8'hf9;
      17'd26944: data = 8'h05;
      17'd26945: data = 8'h0c;
      17'd26946: data = 8'h16;
      17'd26947: data = 8'h16;
      17'd26948: data = 8'h12;
      17'd26949: data = 8'h13;
      17'd26950: data = 8'h0c;
      17'd26951: data = 8'h01;
      17'd26952: data = 8'h02;
      17'd26953: data = 8'h05;
      17'd26954: data = 8'h04;
      17'd26955: data = 8'h04;
      17'd26956: data = 8'hfe;
      17'd26957: data = 8'h01;
      17'd26958: data = 8'h05;
      17'd26959: data = 8'h04;
      17'd26960: data = 8'h0c;
      17'd26961: data = 8'h0e;
      17'd26962: data = 8'h0c;
      17'd26963: data = 8'h06;
      17'd26964: data = 8'h02;
      17'd26965: data = 8'hf9;
      17'd26966: data = 8'hf1;
      17'd26967: data = 8'he9;
      17'd26968: data = 8'he5;
      17'd26969: data = 8'he7;
      17'd26970: data = 8'he7;
      17'd26971: data = 8'hed;
      17'd26972: data = 8'hf9;
      17'd26973: data = 8'hfe;
      17'd26974: data = 8'h01;
      17'd26975: data = 8'h04;
      17'd26976: data = 8'h02;
      17'd26977: data = 8'hfe;
      17'd26978: data = 8'hfe;
      17'd26979: data = 8'hfd;
      17'd26980: data = 8'hf6;
      17'd26981: data = 8'hf9;
      17'd26982: data = 8'hfa;
      17'd26983: data = 8'hf9;
      17'd26984: data = 8'h00;
      17'd26985: data = 8'hfd;
      17'd26986: data = 8'hfa;
      17'd26987: data = 8'h00;
      17'd26988: data = 8'hfe;
      17'd26989: data = 8'h00;
      17'd26990: data = 8'h09;
      17'd26991: data = 8'h05;
      17'd26992: data = 8'h02;
      17'd26993: data = 8'h04;
      17'd26994: data = 8'h05;
      17'd26995: data = 8'h05;
      17'd26996: data = 8'hfe;
      17'd26997: data = 8'h01;
      17'd26998: data = 8'h06;
      17'd26999: data = 8'h0e;
      17'd27000: data = 8'h1b;
      17'd27001: data = 8'h1a;
      17'd27002: data = 8'h1a;
      17'd27003: data = 8'h1c;
      17'd27004: data = 8'h13;
      17'd27005: data = 8'h0e;
      17'd27006: data = 8'h0e;
      17'd27007: data = 8'hfc;
      17'd27008: data = 8'hfa;
      17'd27009: data = 8'h04;
      17'd27010: data = 8'h0a;
      17'd27011: data = 8'h04;
      17'd27012: data = 8'h04;
      17'd27013: data = 8'h1e;
      17'd27014: data = 8'h06;
      17'd27015: data = 8'h00;
      17'd27016: data = 8'h16;
      17'd27017: data = 8'hf6;
      17'd27018: data = 8'hf5;
      17'd27019: data = 8'h0d;
      17'd27020: data = 8'hed;
      17'd27021: data = 8'hfa;
      17'd27022: data = 8'h06;
      17'd27023: data = 8'he4;
      17'd27024: data = 8'h01;
      17'd27025: data = 8'hfd;
      17'd27026: data = 8'hd1;
      17'd27027: data = 8'he5;
      17'd27028: data = 8'hde;
      17'd27029: data = 8'hc4;
      17'd27030: data = 8'hda;
      17'd27031: data = 8'hcb;
      17'd27032: data = 8'hec;
      17'd27033: data = 8'h16;
      17'd27034: data = 8'h0d;
      17'd27035: data = 8'h42;
      17'd27036: data = 8'h54;
      17'd27037: data = 8'h39;
      17'd27038: data = 8'h47;
      17'd27039: data = 8'h3c;
      17'd27040: data = 8'h22;
      17'd27041: data = 8'h2d;
      17'd27042: data = 8'h1b;
      17'd27043: data = 8'h2b;
      17'd27044: data = 8'h2f;
      17'd27045: data = 8'h11;
      17'd27046: data = 8'h27;
      17'd27047: data = 8'h34;
      17'd27048: data = 8'h2b;
      17'd27049: data = 8'h45;
      17'd27050: data = 8'h4f;
      17'd27051: data = 8'h46;
      17'd27052: data = 8'h4a;
      17'd27053: data = 8'h33;
      17'd27054: data = 8'h23;
      17'd27055: data = 8'h15;
      17'd27056: data = 8'hf5;
      17'd27057: data = 8'heb;
      17'd27058: data = 8'hdb;
      17'd27059: data = 8'hc6;
      17'd27060: data = 8'hbd;
      17'd27061: data = 8'hc4;
      17'd27062: data = 8'hd1;
      17'd27063: data = 8'hdb;
      17'd27064: data = 8'he4;
      17'd27065: data = 8'he7;
      17'd27066: data = 8'he3;
      17'd27067: data = 8'hce;
      17'd27068: data = 8'hc5;
      17'd27069: data = 8'hc2;
      17'd27070: data = 8'hb9;
      17'd27071: data = 8'hb5;
      17'd27072: data = 8'hb9;
      17'd27073: data = 8'hb3;
      17'd27074: data = 8'hb0;
      17'd27075: data = 8'hb8;
      17'd27076: data = 8'hc0;
      17'd27077: data = 8'hde;
      17'd27078: data = 8'hf4;
      17'd27079: data = 8'h06;
      17'd27080: data = 8'h22;
      17'd27081: data = 8'h23;
      17'd27082: data = 8'h1c;
      17'd27083: data = 8'h1f;
      17'd27084: data = 8'h15;
      17'd27085: data = 8'h15;
      17'd27086: data = 8'h16;
      17'd27087: data = 8'h16;
      17'd27088: data = 8'h22;
      17'd27089: data = 8'h23;
      17'd27090: data = 8'h2b;
      17'd27091: data = 8'h43;
      17'd27092: data = 8'h4e;
      17'd27093: data = 8'h57;
      17'd27094: data = 8'h60;
      17'd27095: data = 8'h5b;
      17'd27096: data = 8'h54;
      17'd27097: data = 8'h47;
      17'd27098: data = 8'h3a;
      17'd27099: data = 8'h35;
      17'd27100: data = 8'h24;
      17'd27101: data = 8'h13;
      17'd27102: data = 8'h0a;
      17'd27103: data = 8'hf6;
      17'd27104: data = 8'hf1;
      17'd27105: data = 8'hf9;
      17'd27106: data = 8'hfe;
      17'd27107: data = 8'h0a;
      17'd27108: data = 8'h12;
      17'd27109: data = 8'h0d;
      17'd27110: data = 8'h04;
      17'd27111: data = 8'hf5;
      17'd27112: data = 8'he4;
      17'd27113: data = 8'hdb;
      17'd27114: data = 8'hd2;
      17'd27115: data = 8'hc9;
      17'd27116: data = 8'hc4;
      17'd27117: data = 8'hc1;
      17'd27118: data = 8'hc0;
      17'd27119: data = 8'hc6;
      17'd27120: data = 8'hd3;
      17'd27121: data = 8'he2;
      17'd27122: data = 8'hec;
      17'd27123: data = 8'hf5;
      17'd27124: data = 8'hfc;
      17'd27125: data = 8'hfc;
      17'd27126: data = 8'hfc;
      17'd27127: data = 8'h00;
      17'd27128: data = 8'h01;
      17'd27129: data = 8'hfc;
      17'd27130: data = 8'hf6;
      17'd27131: data = 8'hf6;
      17'd27132: data = 8'hf5;
      17'd27133: data = 8'hfc;
      17'd27134: data = 8'h0a;
      17'd27135: data = 8'h1b;
      17'd27136: data = 8'h2b;
      17'd27137: data = 8'h31;
      17'd27138: data = 8'h34;
      17'd27139: data = 8'h33;
      17'd27140: data = 8'h27;
      17'd27141: data = 8'h22;
      17'd27142: data = 8'h1b;
      17'd27143: data = 8'h13;
      17'd27144: data = 8'h0c;
      17'd27145: data = 8'h04;
      17'd27146: data = 8'hfc;
      17'd27147: data = 8'hf6;
      17'd27148: data = 8'hf4;
      17'd27149: data = 8'hf5;
      17'd27150: data = 8'hfa;
      17'd27151: data = 8'hfd;
      17'd27152: data = 8'hfd;
      17'd27153: data = 8'hfa;
      17'd27154: data = 8'hf4;
      17'd27155: data = 8'heb;
      17'd27156: data = 8'hde;
      17'd27157: data = 8'hd8;
      17'd27158: data = 8'hd2;
      17'd27159: data = 8'hc0;
      17'd27160: data = 8'hb4;
      17'd27161: data = 8'hb5;
      17'd27162: data = 8'hc0;
      17'd27163: data = 8'hca;
      17'd27164: data = 8'hda;
      17'd27165: data = 8'hed;
      17'd27166: data = 8'hf6;
      17'd27167: data = 8'hf4;
      17'd27168: data = 8'hf2;
      17'd27169: data = 8'heb;
      17'd27170: data = 8'he5;
      17'd27171: data = 8'he4;
      17'd27172: data = 8'he5;
      17'd27173: data = 8'hed;
      17'd27174: data = 8'heb;
      17'd27175: data = 8'hed;
      17'd27176: data = 8'hfe;
      17'd27177: data = 8'h05;
      17'd27178: data = 8'h05;
      17'd27179: data = 8'h12;
      17'd27180: data = 8'h19;
      17'd27181: data = 8'h1a;
      17'd27182: data = 8'h22;
      17'd27183: data = 8'h1e;
      17'd27184: data = 8'h1c;
      17'd27185: data = 8'h12;
      17'd27186: data = 8'h04;
      17'd27187: data = 8'h04;
      17'd27188: data = 8'hf9;
      17'd27189: data = 8'hf5;
      17'd27190: data = 8'hf9;
      17'd27191: data = 8'hfc;
      17'd27192: data = 8'h00;
      17'd27193: data = 8'h00;
      17'd27194: data = 8'h01;
      17'd27195: data = 8'h01;
      17'd27196: data = 8'hf9;
      17'd27197: data = 8'hf4;
      17'd27198: data = 8'hf1;
      17'd27199: data = 8'hef;
      17'd27200: data = 8'hec;
      17'd27201: data = 8'he9;
      17'd27202: data = 8'he9;
      17'd27203: data = 8'he7;
      17'd27204: data = 8'he9;
      17'd27205: data = 8'hec;
      17'd27206: data = 8'hed;
      17'd27207: data = 8'hed;
      17'd27208: data = 8'hf2;
      17'd27209: data = 8'hf6;
      17'd27210: data = 8'hfc;
      17'd27211: data = 8'hfd;
      17'd27212: data = 8'hfc;
      17'd27213: data = 8'hfa;
      17'd27214: data = 8'hf5;
      17'd27215: data = 8'hf4;
      17'd27216: data = 8'hf4;
      17'd27217: data = 8'hf5;
      17'd27218: data = 8'h00;
      17'd27219: data = 8'h0c;
      17'd27220: data = 8'h0e;
      17'd27221: data = 8'h11;
      17'd27222: data = 8'h0e;
      17'd27223: data = 8'h0c;
      17'd27224: data = 8'h05;
      17'd27225: data = 8'h00;
      17'd27226: data = 8'hfc;
      17'd27227: data = 8'hfa;
      17'd27228: data = 8'h02;
      17'd27229: data = 8'h04;
      17'd27230: data = 8'h01;
      17'd27231: data = 8'h0c;
      17'd27232: data = 8'h06;
      17'd27233: data = 8'h05;
      17'd27234: data = 8'h0a;
      17'd27235: data = 8'h01;
      17'd27236: data = 8'h12;
      17'd27237: data = 8'h15;
      17'd27238: data = 8'h0c;
      17'd27239: data = 8'h19;
      17'd27240: data = 8'h02;
      17'd27241: data = 8'hf6;
      17'd27242: data = 8'h11;
      17'd27243: data = 8'hf9;
      17'd27244: data = 8'hf4;
      17'd27245: data = 8'h16;
      17'd27246: data = 8'hf6;
      17'd27247: data = 8'h01;
      17'd27248: data = 8'h23;
      17'd27249: data = 8'h0c;
      17'd27250: data = 8'hfe;
      17'd27251: data = 8'h02;
      17'd27252: data = 8'hfa;
      17'd27253: data = 8'heb;
      17'd27254: data = 8'hef;
      17'd27255: data = 8'hec;
      17'd27256: data = 8'hf5;
      17'd27257: data = 8'h1c;
      17'd27258: data = 8'h13;
      17'd27259: data = 8'h01;
      17'd27260: data = 8'h24;
      17'd27261: data = 8'h05;
      17'd27262: data = 8'hed;
      17'd27263: data = 8'hf9;
      17'd27264: data = 8'hd6;
      17'd27265: data = 8'hd2;
      17'd27266: data = 8'he7;
      17'd27267: data = 8'hc9;
      17'd27268: data = 8'hd5;
      17'd27269: data = 8'hfe;
      17'd27270: data = 8'hf1;
      17'd27271: data = 8'h26;
      17'd27272: data = 8'h4f;
      17'd27273: data = 8'h47;
      17'd27274: data = 8'h60;
      17'd27275: data = 8'h57;
      17'd27276: data = 8'h39;
      17'd27277: data = 8'h42;
      17'd27278: data = 8'h24;
      17'd27279: data = 8'h23;
      17'd27280: data = 8'h1e;
      17'd27281: data = 8'h0e;
      17'd27282: data = 8'h16;
      17'd27283: data = 8'h13;
      17'd27284: data = 8'h24;
      17'd27285: data = 8'h34;
      17'd27286: data = 8'h4a;
      17'd27287: data = 8'h54;
      17'd27288: data = 8'h57;
      17'd27289: data = 8'h43;
      17'd27290: data = 8'h39;
      17'd27291: data = 8'h24;
      17'd27292: data = 8'h01;
      17'd27293: data = 8'hf6;
      17'd27294: data = 8'he3;
      17'd27295: data = 8'hcd;
      17'd27296: data = 8'hc2;
      17'd27297: data = 8'hb3;
      17'd27298: data = 8'hb4;
      17'd27299: data = 8'hc4;
      17'd27300: data = 8'hd5;
      17'd27301: data = 8'he5;
      17'd27302: data = 8'hf2;
      17'd27303: data = 8'hed;
      17'd27304: data = 8'he2;
      17'd27305: data = 8'hd6;
      17'd27306: data = 8'hc6;
      17'd27307: data = 8'hbd;
      17'd27308: data = 8'hb5;
      17'd27309: data = 8'hb0;
      17'd27310: data = 8'ha8;
      17'd27311: data = 8'hac;
      17'd27312: data = 8'hae;
      17'd27313: data = 8'hbc;
      17'd27314: data = 8'hd8;
      17'd27315: data = 8'hf2;
      17'd27316: data = 8'h0d;
      17'd27317: data = 8'h1e;
      17'd27318: data = 8'h29;
      17'd27319: data = 8'h24;
      17'd27320: data = 8'h1b;
      17'd27321: data = 8'h23;
      17'd27322: data = 8'h1b;
      17'd27323: data = 8'h19;
      17'd27324: data = 8'h1c;
      17'd27325: data = 8'h12;
      17'd27326: data = 8'h15;
      17'd27327: data = 8'h22;
      17'd27328: data = 8'h2b;
      17'd27329: data = 8'h43;
      17'd27330: data = 8'h54;
      17'd27331: data = 8'h5a;
      17'd27332: data = 8'h5d;
      17'd27333: data = 8'h57;
      17'd27334: data = 8'h4a;
      17'd27335: data = 8'h40;
      17'd27336: data = 8'h31;
      17'd27337: data = 8'h23;
      17'd27338: data = 8'h15;
      17'd27339: data = 8'h02;
      17'd27340: data = 8'hf5;
      17'd27341: data = 8'hec;
      17'd27342: data = 8'hed;
      17'd27343: data = 8'hf6;
      17'd27344: data = 8'hfe;
      17'd27345: data = 8'h05;
      17'd27346: data = 8'h0c;
      17'd27347: data = 8'h04;
      17'd27348: data = 8'hfa;
      17'd27349: data = 8'hed;
      17'd27350: data = 8'he3;
      17'd27351: data = 8'hda;
      17'd27352: data = 8'hce;
      17'd27353: data = 8'hc9;
      17'd27354: data = 8'hc1;
      17'd27355: data = 8'hbc;
      17'd27356: data = 8'hc1;
      17'd27357: data = 8'hcd;
      17'd27358: data = 8'hdc;
      17'd27359: data = 8'hec;
      17'd27360: data = 8'hf9;
      17'd27361: data = 8'hfa;
      17'd27362: data = 8'hfd;
      17'd27363: data = 8'h00;
      17'd27364: data = 8'h02;
      17'd27365: data = 8'h01;
      17'd27366: data = 8'h01;
      17'd27367: data = 8'hfc;
      17'd27368: data = 8'hf5;
      17'd27369: data = 8'hf4;
      17'd27370: data = 8'hf9;
      17'd27371: data = 8'h02;
      17'd27372: data = 8'h12;
      17'd27373: data = 8'h1e;
      17'd27374: data = 8'h29;
      17'd27375: data = 8'h2f;
      17'd27376: data = 8'h2d;
      17'd27377: data = 8'h29;
      17'd27378: data = 8'h26;
      17'd27379: data = 8'h1f;
      17'd27380: data = 8'h16;
      17'd27381: data = 8'h0e;
      17'd27382: data = 8'h02;
      17'd27383: data = 8'hfa;
      17'd27384: data = 8'hf2;
      17'd27385: data = 8'hf1;
      17'd27386: data = 8'hef;
      17'd27387: data = 8'hef;
      17'd27388: data = 8'hf5;
      17'd27389: data = 8'hf1;
      17'd27390: data = 8'hec;
      17'd27391: data = 8'heb;
      17'd27392: data = 8'hec;
      17'd27393: data = 8'he5;
      17'd27394: data = 8'he3;
      17'd27395: data = 8'hdb;
      17'd27396: data = 8'hd1;
      17'd27397: data = 8'hc4;
      17'd27398: data = 8'hbc;
      17'd27399: data = 8'hbd;
      17'd27400: data = 8'hc6;
      17'd27401: data = 8'hcd;
      17'd27402: data = 8'hd6;
      17'd27403: data = 8'hdb;
      17'd27404: data = 8'he2;
      17'd27405: data = 8'hec;
      17'd27406: data = 8'hf2;
      17'd27407: data = 8'hfd;
      17'd27408: data = 8'h04;
      17'd27409: data = 8'h00;
      17'd27410: data = 8'h02;
      17'd27411: data = 8'h01;
      17'd27412: data = 8'hfc;
      17'd27413: data = 8'hfc;
      17'd27414: data = 8'hfa;
      17'd27415: data = 8'hfd;
      17'd27416: data = 8'h01;
      17'd27417: data = 8'h0a;
      17'd27418: data = 8'h12;
      17'd27419: data = 8'h19;
      17'd27420: data = 8'h1c;
      17'd27421: data = 8'h1e;
      17'd27422: data = 8'h1b;
      17'd27423: data = 8'h13;
      17'd27424: data = 8'h0d;
      17'd27425: data = 8'h05;
      17'd27426: data = 8'hfe;
      17'd27427: data = 8'hf9;
      17'd27428: data = 8'hf2;
      17'd27429: data = 8'hec;
      17'd27430: data = 8'hec;
      17'd27431: data = 8'hec;
      17'd27432: data = 8'hed;
      17'd27433: data = 8'hef;
      17'd27434: data = 8'hf6;
      17'd27435: data = 8'hfc;
      17'd27436: data = 8'hfc;
      17'd27437: data = 8'hfa;
      17'd27438: data = 8'hf2;
      17'd27439: data = 8'hef;
      17'd27440: data = 8'hec;
      17'd27441: data = 8'he4;
      17'd27442: data = 8'he3;
      17'd27443: data = 8'he2;
      17'd27444: data = 8'he4;
      17'd27445: data = 8'he7;
      17'd27446: data = 8'hf1;
      17'd27447: data = 8'hf6;
      17'd27448: data = 8'hfa;
      17'd27449: data = 8'h05;
      17'd27450: data = 8'h04;
      17'd27451: data = 8'h02;
      17'd27452: data = 8'h05;
      17'd27453: data = 8'h02;
      17'd27454: data = 8'h00;
      17'd27455: data = 8'hfe;
      17'd27456: data = 8'h00;
      17'd27457: data = 8'hfd;
      17'd27458: data = 8'hfc;
      17'd27459: data = 8'hfa;
      17'd27460: data = 8'hfd;
      17'd27461: data = 8'h00;
      17'd27462: data = 8'h00;
      17'd27463: data = 8'h0a;
      17'd27464: data = 8'h0e;
      17'd27465: data = 8'h11;
      17'd27466: data = 8'h19;
      17'd27467: data = 8'h11;
      17'd27468: data = 8'h0c;
      17'd27469: data = 8'h06;
      17'd27470: data = 8'h00;
      17'd27471: data = 8'hfc;
      17'd27472: data = 8'hf6;
      17'd27473: data = 8'h01;
      17'd27474: data = 8'h05;
      17'd27475: data = 8'h05;
      17'd27476: data = 8'h12;
      17'd27477: data = 8'h0a;
      17'd27478: data = 8'h0d;
      17'd27479: data = 8'h0c;
      17'd27480: data = 8'hfe;
      17'd27481: data = 8'h16;
      17'd27482: data = 8'h12;
      17'd27483: data = 8'h01;
      17'd27484: data = 8'h0c;
      17'd27485: data = 8'hfe;
      17'd27486: data = 8'hf9;
      17'd27487: data = 8'hf2;
      17'd27488: data = 8'hec;
      17'd27489: data = 8'hfd;
      17'd27490: data = 8'hfc;
      17'd27491: data = 8'hfc;
      17'd27492: data = 8'h0a;
      17'd27493: data = 8'h16;
      17'd27494: data = 8'h11;
      17'd27495: data = 8'h02;
      17'd27496: data = 8'h0a;
      17'd27497: data = 8'h11;
      17'd27498: data = 8'hfa;
      17'd27499: data = 8'hdb;
      17'd27500: data = 8'hd1;
      17'd27501: data = 8'hc9;
      17'd27502: data = 8'hbb;
      17'd27503: data = 8'hb0;
      17'd27504: data = 8'hd1;
      17'd27505: data = 8'h05;
      17'd27506: data = 8'h1f;
      17'd27507: data = 8'h40;
      17'd27508: data = 8'h67;
      17'd27509: data = 8'h5c;
      17'd27510: data = 8'h57;
      17'd27511: data = 8'h4a;
      17'd27512: data = 8'h36;
      17'd27513: data = 8'h33;
      17'd27514: data = 8'h13;
      17'd27515: data = 8'h12;
      17'd27516: data = 8'h13;
      17'd27517: data = 8'h13;
      17'd27518: data = 8'h19;
      17'd27519: data = 8'h26;
      17'd27520: data = 8'h3a;
      17'd27521: data = 8'h46;
      17'd27522: data = 8'h5a;
      17'd27523: data = 8'h63;
      17'd27524: data = 8'h5a;
      17'd27525: data = 8'h4e;
      17'd27526: data = 8'h47;
      17'd27527: data = 8'h2c;
      17'd27528: data = 8'h09;
      17'd27529: data = 8'he4;
      17'd27530: data = 8'hcb;
      17'd27531: data = 8'hb3;
      17'd27532: data = 8'h9f;
      17'd27533: data = 8'hb1;
      17'd27534: data = 8'hca;
      17'd27535: data = 8'hda;
      17'd27536: data = 8'he7;
      17'd27537: data = 8'hf4;
      17'd27538: data = 8'hef;
      17'd27539: data = 8'hdc;
      17'd27540: data = 8'hd2;
      17'd27541: data = 8'hcb;
      17'd27542: data = 8'hc0;
      17'd27543: data = 8'hac;
      17'd27544: data = 8'ha8;
      17'd27545: data = 8'h9f;
      17'd27546: data = 8'h92;
      17'd27547: data = 8'h95;
      17'd27548: data = 8'ha3;
      17'd27549: data = 8'hbc;
      17'd27550: data = 8'hd3;
      17'd27551: data = 8'hf1;
      17'd27552: data = 8'h0e;
      17'd27553: data = 8'h1a;
      17'd27554: data = 8'h1f;
      17'd27555: data = 8'h27;
      17'd27556: data = 8'h23;
      17'd27557: data = 8'h1b;
      17'd27558: data = 8'h12;
      17'd27559: data = 8'h0d;
      17'd27560: data = 8'h0c;
      17'd27561: data = 8'h0a;
      17'd27562: data = 8'h1b;
      17'd27563: data = 8'h2c;
      17'd27564: data = 8'h3d;
      17'd27565: data = 8'h4f;
      17'd27566: data = 8'h5c;
      17'd27567: data = 8'h64;
      17'd27568: data = 8'h63;
      17'd27569: data = 8'h65;
      17'd27570: data = 8'h63;
      17'd27571: data = 8'h52;
      17'd27572: data = 8'h3d;
      17'd27573: data = 8'h2c;
      17'd27574: data = 8'h13;
      17'd27575: data = 8'hfe;
      17'd27576: data = 8'hfa;
      17'd27577: data = 8'hf6;
      17'd27578: data = 8'hfa;
      17'd27579: data = 8'h04;
      17'd27580: data = 8'h0d;
      17'd27581: data = 8'h11;
      17'd27582: data = 8'h0a;
      17'd27583: data = 8'h0a;
      17'd27584: data = 8'h02;
      17'd27585: data = 8'hf4;
      17'd27586: data = 8'he4;
      17'd27587: data = 8'hd5;
      17'd27588: data = 8'hc4;
      17'd27589: data = 8'hb5;
      17'd27590: data = 8'hb3;
      17'd27591: data = 8'hb8;
      17'd27592: data = 8'hc0;
      17'd27593: data = 8'hc2;
      17'd27594: data = 8'hce;
      17'd27595: data = 8'hdb;
      17'd27596: data = 8'he4;
      17'd27597: data = 8'hf1;
      17'd27598: data = 8'hfd;
      17'd27599: data = 8'h04;
      17'd27600: data = 8'h00;
      17'd27601: data = 8'hfe;
      17'd27602: data = 8'hfa;
      17'd27603: data = 8'hec;
      17'd27604: data = 8'he7;
      17'd27605: data = 8'hec;
      17'd27606: data = 8'hf2;
      17'd27607: data = 8'h01;
      17'd27608: data = 8'h11;
      17'd27609: data = 8'h24;
      17'd27610: data = 8'h2d;
      17'd27611: data = 8'h35;
      17'd27612: data = 8'h3d;
      17'd27613: data = 8'h3c;
      17'd27614: data = 8'h35;
      17'd27615: data = 8'h2c;
      17'd27616: data = 8'h26;
      17'd27617: data = 8'h1b;
      17'd27618: data = 8'h0e;
      17'd27619: data = 8'h00;
      17'd27620: data = 8'hf4;
      17'd27621: data = 8'hf4;
      17'd27622: data = 8'hf1;
      17'd27623: data = 8'heb;
      17'd27624: data = 8'hf1;
      17'd27625: data = 8'hfc;
      17'd27626: data = 8'hfd;
      17'd27627: data = 8'hfa;
      17'd27628: data = 8'hf9;
      17'd27629: data = 8'hf4;
      17'd27630: data = 8'he4;
      17'd27631: data = 8'hd5;
      17'd27632: data = 8'hc9;
      17'd27633: data = 8'hbb;
      17'd27634: data = 8'hb1;
      17'd27635: data = 8'hb4;
      17'd27636: data = 8'hb8;
      17'd27637: data = 8'hbc;
      17'd27638: data = 8'hc9;
      17'd27639: data = 8'hd1;
      17'd27640: data = 8'hdc;
      17'd27641: data = 8'he5;
      17'd27642: data = 8'he7;
      17'd27643: data = 8'hf2;
      17'd27644: data = 8'hf2;
      17'd27645: data = 8'hed;
      17'd27646: data = 8'hf2;
      17'd27647: data = 8'hef;
      17'd27648: data = 8'he7;
      17'd27649: data = 8'he7;
      17'd27650: data = 8'hf2;
      17'd27651: data = 8'hfa;
      17'd27652: data = 8'h02;
      17'd27653: data = 8'h11;
      17'd27654: data = 8'h1c;
      17'd27655: data = 8'h26;
      17'd27656: data = 8'h24;
      17'd27657: data = 8'h27;
      17'd27658: data = 8'h24;
      17'd27659: data = 8'h19;
      17'd27660: data = 8'h11;
      17'd27661: data = 8'h04;
      17'd27662: data = 8'hfd;
      17'd27663: data = 8'hf5;
      17'd27664: data = 8'hf4;
      17'd27665: data = 8'hf9;
      17'd27666: data = 8'hf5;
      17'd27667: data = 8'hfd;
      17'd27668: data = 8'h05;
      17'd27669: data = 8'h06;
      17'd27670: data = 8'h06;
      17'd27671: data = 8'h04;
      17'd27672: data = 8'h02;
      17'd27673: data = 8'hfd;
      17'd27674: data = 8'hf2;
      17'd27675: data = 8'hed;
      17'd27676: data = 8'he5;
      17'd27677: data = 8'he0;
      17'd27678: data = 8'hde;
      17'd27679: data = 8'hda;
      17'd27680: data = 8'he0;
      17'd27681: data = 8'he5;
      17'd27682: data = 8'hec;
      17'd27683: data = 8'hf5;
      17'd27684: data = 8'hfc;
      17'd27685: data = 8'hfe;
      17'd27686: data = 8'h01;
      17'd27687: data = 8'hfa;
      17'd27688: data = 8'hf6;
      17'd27689: data = 8'hfa;
      17'd27690: data = 8'hf1;
      17'd27691: data = 8'hf1;
      17'd27692: data = 8'hed;
      17'd27693: data = 8'hec;
      17'd27694: data = 8'hf2;
      17'd27695: data = 8'hf2;
      17'd27696: data = 8'h01;
      17'd27697: data = 8'h09;
      17'd27698: data = 8'h0a;
      17'd27699: data = 8'h1a;
      17'd27700: data = 8'h15;
      17'd27701: data = 8'h12;
      17'd27702: data = 8'h16;
      17'd27703: data = 8'h05;
      17'd27704: data = 8'h0a;
      17'd27705: data = 8'h02;
      17'd27706: data = 8'h00;
      17'd27707: data = 8'h16;
      17'd27708: data = 8'h06;
      17'd27709: data = 8'h0c;
      17'd27710: data = 8'h15;
      17'd27711: data = 8'h01;
      17'd27712: data = 8'h19;
      17'd27713: data = 8'h22;
      17'd27714: data = 8'h11;
      17'd27715: data = 8'h1e;
      17'd27716: data = 8'h11;
      17'd27717: data = 8'hfd;
      17'd27718: data = 8'h15;
      17'd27719: data = 8'hfc;
      17'd27720: data = 8'heb;
      17'd27721: data = 8'h1e;
      17'd27722: data = 8'h01;
      17'd27723: data = 8'hf6;
      17'd27724: data = 8'h16;
      17'd27725: data = 8'hf5;
      17'd27726: data = 8'hfe;
      17'd27727: data = 8'h02;
      17'd27728: data = 8'he0;
      17'd27729: data = 8'h04;
      17'd27730: data = 8'hfd;
      17'd27731: data = 8'he9;
      17'd27732: data = 8'h22;
      17'd27733: data = 8'h06;
      17'd27734: data = 8'hdc;
      17'd27735: data = 8'hf2;
      17'd27736: data = 8'hd8;
      17'd27737: data = 8'hb9;
      17'd27738: data = 8'hce;
      17'd27739: data = 8'hc2;
      17'd27740: data = 8'he0;
      17'd27741: data = 8'h0d;
      17'd27742: data = 8'h0e;
      17'd27743: data = 8'h47;
      17'd27744: data = 8'h5c;
      17'd27745: data = 8'h3a;
      17'd27746: data = 8'h4a;
      17'd27747: data = 8'h3a;
      17'd27748: data = 8'h1e;
      17'd27749: data = 8'h27;
      17'd27750: data = 8'h26;
      17'd27751: data = 8'h2c;
      17'd27752: data = 8'h34;
      17'd27753: data = 8'h23;
      17'd27754: data = 8'h26;
      17'd27755: data = 8'h36;
      17'd27756: data = 8'h26;
      17'd27757: data = 8'h3e;
      17'd27758: data = 8'h52;
      17'd27759: data = 8'h4e;
      17'd27760: data = 8'h5c;
      17'd27761: data = 8'h57;
      17'd27762: data = 8'h43;
      17'd27763: data = 8'h31;
      17'd27764: data = 8'h05;
      17'd27765: data = 8'hfc;
      17'd27766: data = 8'he5;
      17'd27767: data = 8'hc2;
      17'd27768: data = 8'hce;
      17'd27769: data = 8'hd2;
      17'd27770: data = 8'hcb;
      17'd27771: data = 8'he2;
      17'd27772: data = 8'he4;
      17'd27773: data = 8'he3;
      17'd27774: data = 8'hdc;
      17'd27775: data = 8'hca;
      17'd27776: data = 8'hcd;
      17'd27777: data = 8'hc4;
      17'd27778: data = 8'hb1;
      17'd27779: data = 8'hb8;
      17'd27780: data = 8'hb0;
      17'd27781: data = 8'h99;
      17'd27782: data = 8'h9b;
      17'd27783: data = 8'h94;
      17'd27784: data = 8'h92;
      17'd27785: data = 8'ha4;
      17'd27786: data = 8'hbb;
      17'd27787: data = 8'hda;
      17'd27788: data = 8'hf2;
      17'd27789: data = 8'hf9;
      17'd27790: data = 8'h0e;
      17'd27791: data = 8'h0e;
      17'd27792: data = 8'h01;
      17'd27793: data = 8'h0e;
      17'd27794: data = 8'h0e;
      17'd27795: data = 8'h09;
      17'd27796: data = 8'h0e;
      17'd27797: data = 8'h1b;
      17'd27798: data = 8'h24;
      17'd27799: data = 8'h31;
      17'd27800: data = 8'h3e;
      17'd27801: data = 8'h52;
      17'd27802: data = 8'h56;
      17'd27803: data = 8'h5a;
      17'd27804: data = 8'h67;
      17'd27805: data = 8'h6c;
      17'd27806: data = 8'h68;
      17'd27807: data = 8'h68;
      17'd27808: data = 8'h5d;
      17'd27809: data = 8'h4f;
      17'd27810: data = 8'h3a;
      17'd27811: data = 8'h27;
      17'd27812: data = 8'h23;
      17'd27813: data = 8'h12;
      17'd27814: data = 8'h16;
      17'd27815: data = 8'h24;
      17'd27816: data = 8'h22;
      17'd27817: data = 8'h1f;
      17'd27818: data = 8'h1e;
      17'd27819: data = 8'h12;
      17'd27820: data = 8'h05;
      17'd27821: data = 8'hf9;
      17'd27822: data = 8'hec;
      17'd27823: data = 8'hde;
      17'd27824: data = 8'hcd;
      17'd27825: data = 8'hc5;
      17'd27826: data = 8'hc0;
      17'd27827: data = 8'hb1;
      17'd27828: data = 8'hb3;
      17'd27829: data = 8'hb9;
      17'd27830: data = 8'hb4;
      17'd27831: data = 8'hbd;
      17'd27832: data = 8'hc1;
      17'd27833: data = 8'hcb;
      17'd27834: data = 8'hda;
      17'd27835: data = 8'hde;
      17'd27836: data = 8'he4;
      17'd27837: data = 8'he4;
      17'd27838: data = 8'hdc;
      17'd27839: data = 8'hd8;
      17'd27840: data = 8'hd8;
      17'd27841: data = 8'hdb;
      17'd27842: data = 8'he4;
      17'd27843: data = 8'hf4;
      17'd27844: data = 8'h02;
      17'd27845: data = 8'h12;
      17'd27846: data = 8'h1c;
      17'd27847: data = 8'h26;
      17'd27848: data = 8'h2f;
      17'd27849: data = 8'h33;
      17'd27850: data = 8'h34;
      17'd27851: data = 8'h3a;
      17'd27852: data = 8'h39;
      17'd27853: data = 8'h33;
      17'd27854: data = 8'h2b;
      17'd27855: data = 8'h1f;
      17'd27856: data = 8'h16;
      17'd27857: data = 8'h11;
      17'd27858: data = 8'h15;
      17'd27859: data = 8'h15;
      17'd27860: data = 8'h13;
      17'd27861: data = 8'h19;
      17'd27862: data = 8'h1b;
      17'd27863: data = 8'h15;
      17'd27864: data = 8'h0e;
      17'd27865: data = 8'h04;
      17'd27866: data = 8'hf6;
      17'd27867: data = 8'heb;
      17'd27868: data = 8'hdc;
      17'd27869: data = 8'hd2;
      17'd27870: data = 8'hc6;
      17'd27871: data = 8'hbd;
      17'd27872: data = 8'hb9;
      17'd27873: data = 8'hb8;
      17'd27874: data = 8'hb5;
      17'd27875: data = 8'hc0;
      17'd27876: data = 8'hc4;
      17'd27877: data = 8'hce;
      17'd27878: data = 8'hd2;
      17'd27879: data = 8'hce;
      17'd27880: data = 8'hd2;
      17'd27881: data = 8'hc6;
      17'd27882: data = 8'hc2;
      17'd27883: data = 8'hca;
      17'd27884: data = 8'hc6;
      17'd27885: data = 8'hca;
      17'd27886: data = 8'hd6;
      17'd27887: data = 8'hde;
      17'd27888: data = 8'he7;
      17'd27889: data = 8'hf5;
      17'd27890: data = 8'hfc;
      17'd27891: data = 8'h06;
      17'd27892: data = 8'h0e;
      17'd27893: data = 8'h16;
      17'd27894: data = 8'h1e;
      17'd27895: data = 8'h1e;
      17'd27896: data = 8'h19;
      17'd27897: data = 8'h19;
      17'd27898: data = 8'h12;
      17'd27899: data = 8'h09;
      17'd27900: data = 8'h0c;
      17'd27901: data = 8'h12;
      17'd27902: data = 8'h16;
      17'd27903: data = 8'h1b;
      17'd27904: data = 8'h26;
      17'd27905: data = 8'h27;
      17'd27906: data = 8'h29;
      17'd27907: data = 8'h29;
      17'd27908: data = 8'h22;
      17'd27909: data = 8'h19;
      17'd27910: data = 8'h11;
      17'd27911: data = 8'h0a;
      17'd27912: data = 8'h02;
      17'd27913: data = 8'hfe;
      17'd27914: data = 8'hfd;
      17'd27915: data = 8'hfa;
      17'd27916: data = 8'hf5;
      17'd27917: data = 8'hf4;
      17'd27918: data = 8'hf4;
      17'd27919: data = 8'hf5;
      17'd27920: data = 8'hf4;
      17'd27921: data = 8'hf4;
      17'd27922: data = 8'hf4;
      17'd27923: data = 8'hef;
      17'd27924: data = 8'heb;
      17'd27925: data = 8'he5;
      17'd27926: data = 8'he0;
      17'd27927: data = 8'hd8;
      17'd27928: data = 8'hd5;
      17'd27929: data = 8'hd6;
      17'd27930: data = 8'hda;
      17'd27931: data = 8'hde;
      17'd27932: data = 8'he4;
      17'd27933: data = 8'hed;
      17'd27934: data = 8'hf5;
      17'd27935: data = 8'hf6;
      17'd27936: data = 8'hf9;
      17'd27937: data = 8'hfd;
      17'd27938: data = 8'hfe;
      17'd27939: data = 8'hfa;
      17'd27940: data = 8'hfc;
      17'd27941: data = 8'h04;
      17'd27942: data = 8'h05;
      17'd27943: data = 8'h01;
      17'd27944: data = 8'h09;
      17'd27945: data = 8'h0e;
      17'd27946: data = 8'h16;
      17'd27947: data = 8'h15;
      17'd27948: data = 8'h15;
      17'd27949: data = 8'h27;
      17'd27950: data = 8'h1f;
      17'd27951: data = 8'h13;
      17'd27952: data = 8'h22;
      17'd27953: data = 8'h24;
      17'd27954: data = 8'h1c;
      17'd27955: data = 8'h1e;
      17'd27956: data = 8'h1a;
      17'd27957: data = 8'h22;
      17'd27958: data = 8'h1a;
      17'd27959: data = 8'h0e;
      17'd27960: data = 8'h13;
      17'd27961: data = 8'h05;
      17'd27962: data = 8'hfe;
      17'd27963: data = 8'h09;
      17'd27964: data = 8'h05;
      17'd27965: data = 8'h0a;
      17'd27966: data = 8'h12;
      17'd27967: data = 8'h09;
      17'd27968: data = 8'h0c;
      17'd27969: data = 8'h0c;
      17'd27970: data = 8'h05;
      17'd27971: data = 8'hf4;
      17'd27972: data = 8'hda;
      17'd27973: data = 8'hd2;
      17'd27974: data = 8'hd2;
      17'd27975: data = 8'hc5;
      17'd27976: data = 8'hc1;
      17'd27977: data = 8'hd3;
      17'd27978: data = 8'hec;
      17'd27979: data = 8'hf2;
      17'd27980: data = 8'h05;
      17'd27981: data = 8'h24;
      17'd27982: data = 8'h29;
      17'd27983: data = 8'h26;
      17'd27984: data = 8'h2b;
      17'd27985: data = 8'h24;
      17'd27986: data = 8'h1b;
      17'd27987: data = 8'h16;
      17'd27988: data = 8'h12;
      17'd27989: data = 8'h12;
      17'd27990: data = 8'h09;
      17'd27991: data = 8'h0e;
      17'd27992: data = 8'h1a;
      17'd27993: data = 8'h23;
      17'd27994: data = 8'h34;
      17'd27995: data = 8'h46;
      17'd27996: data = 8'h4e;
      17'd27997: data = 8'h53;
      17'd27998: data = 8'h5a;
      17'd27999: data = 8'h5a;
      17'd28000: data = 8'h43;
      17'd28001: data = 8'h2f;
      17'd28002: data = 8'h1c;
      17'd28003: data = 8'h0e;
      17'd28004: data = 8'hfd;
      17'd28005: data = 8'hf1;
      17'd28006: data = 8'hf6;
      17'd28007: data = 8'hf4;
      17'd28008: data = 8'hf1;
      17'd28009: data = 8'hfc;
      17'd28010: data = 8'hfe;
      17'd28011: data = 8'hfc;
      17'd28012: data = 8'hfe;
      17'd28013: data = 8'hf5;
      17'd28014: data = 8'hed;
      17'd28015: data = 8'he0;
      17'd28016: data = 8'hd5;
      17'd28017: data = 8'hc6;
      17'd28018: data = 8'hb8;
      17'd28019: data = 8'ha4;
      17'd28020: data = 8'ha1;
      17'd28021: data = 8'ha1;
      17'd28022: data = 8'ha6;
      17'd28023: data = 8'hb0;
      17'd28024: data = 8'hbd;
      17'd28025: data = 8'hcb;
      17'd28026: data = 8'hd8;
      17'd28027: data = 8'he2;
      17'd28028: data = 8'he7;
      17'd28029: data = 8'he7;
      17'd28030: data = 8'he4;
      17'd28031: data = 8'he3;
      17'd28032: data = 8'he3;
      17'd28033: data = 8'he7;
      17'd28034: data = 8'hf1;
      17'd28035: data = 8'hf9;
      17'd28036: data = 8'heb;
      17'd28037: data = 8'heb;
      17'd28038: data = 8'hf9;
      17'd28039: data = 8'h15;
      17'd28040: data = 8'h34;
      17'd28041: data = 8'h4e;
      17'd28042: data = 8'h5d;
      17'd28043: data = 8'h72;
      17'd28044: data = 8'h6d;
      17'd28045: data = 8'h4b;
      17'd28046: data = 8'h40;
      17'd28047: data = 8'h42;
      17'd28048: data = 8'h31;
      17'd28049: data = 8'h31;
      17'd28050: data = 8'h39;
      17'd28051: data = 8'h29;
      17'd28052: data = 8'h31;
      17'd28053: data = 8'h46;
      17'd28054: data = 8'h3d;
      17'd28055: data = 8'h3c;
      17'd28056: data = 8'h4e;
      17'd28057: data = 8'h42;
      17'd28058: data = 8'h2d;
      17'd28059: data = 8'h2f;
      17'd28060: data = 8'h2d;
      17'd28061: data = 8'h1a;
      17'd28062: data = 8'h04;
      17'd28063: data = 8'hfc;
      17'd28064: data = 8'heb;
      17'd28065: data = 8'hcb;
      17'd28066: data = 8'hc4;
      17'd28067: data = 8'hc4;
      17'd28068: data = 8'hcd;
      17'd28069: data = 8'hdb;
      17'd28070: data = 8'hdc;
      17'd28071: data = 8'hd6;
      17'd28072: data = 8'hd6;
      17'd28073: data = 8'hd3;
      17'd28074: data = 8'hca;
      17'd28075: data = 8'hc1;
      17'd28076: data = 8'hc0;
      17'd28077: data = 8'hc2;
      17'd28078: data = 8'hbd;
      17'd28079: data = 8'hb9;
      17'd28080: data = 8'hb3;
      17'd28081: data = 8'hb9;
      17'd28082: data = 8'hc1;
      17'd28083: data = 8'hc6;
      17'd28084: data = 8'hd3;
      17'd28085: data = 8'he7;
      17'd28086: data = 8'hf4;
      17'd28087: data = 8'h00;
      17'd28088: data = 8'h06;
      17'd28089: data = 8'h11;
      17'd28090: data = 8'h13;
      17'd28091: data = 8'h0a;
      17'd28092: data = 8'h09;
      17'd28093: data = 8'h09;
      17'd28094: data = 8'h02;
      17'd28095: data = 8'h02;
      17'd28096: data = 8'h0d;
      17'd28097: data = 8'h16;
      17'd28098: data = 8'h1f;
      17'd28099: data = 8'h29;
      17'd28100: data = 8'h31;
      17'd28101: data = 8'h33;
      17'd28102: data = 8'h33;
      17'd28103: data = 8'h33;
      17'd28104: data = 8'h31;
      17'd28105: data = 8'h26;
      17'd28106: data = 8'h1c;
      17'd28107: data = 8'h15;
      17'd28108: data = 8'h09;
      17'd28109: data = 8'hfd;
      17'd28110: data = 8'hf5;
      17'd28111: data = 8'hf1;
      17'd28112: data = 8'hef;
      17'd28113: data = 8'hef;
      17'd28114: data = 8'hf9;
      17'd28115: data = 8'hfa;
      17'd28116: data = 8'hf5;
      17'd28117: data = 8'hf6;
      17'd28118: data = 8'hef;
      17'd28119: data = 8'he4;
      17'd28120: data = 8'hdb;
      17'd28121: data = 8'hd3;
      17'd28122: data = 8'hca;
      17'd28123: data = 8'hc0;
      17'd28124: data = 8'hbd;
      17'd28125: data = 8'hc0;
      17'd28126: data = 8'hc4;
      17'd28127: data = 8'hc5;
      17'd28128: data = 8'hce;
      17'd28129: data = 8'hd5;
      17'd28130: data = 8'hd5;
      17'd28131: data = 8'hdc;
      17'd28132: data = 8'hde;
      17'd28133: data = 8'hdc;
      17'd28134: data = 8'hdc;
      17'd28135: data = 8'hdc;
      17'd28136: data = 8'hda;
      17'd28137: data = 8'hda;
      17'd28138: data = 8'hdc;
      17'd28139: data = 8'he0;
      17'd28140: data = 8'he5;
      17'd28141: data = 8'hef;
      17'd28142: data = 8'hfa;
      17'd28143: data = 8'h05;
      17'd28144: data = 8'h0d;
      17'd28145: data = 8'h13;
      17'd28146: data = 8'h1a;
      17'd28147: data = 8'h19;
      17'd28148: data = 8'h1a;
      17'd28149: data = 8'h1a;
      17'd28150: data = 8'h15;
      17'd28151: data = 8'h16;
      17'd28152: data = 8'h16;
      17'd28153: data = 8'h16;
      17'd28154: data = 8'h19;
      17'd28155: data = 8'h19;
      17'd28156: data = 8'h19;
      17'd28157: data = 8'h1c;
      17'd28158: data = 8'h22;
      17'd28159: data = 8'h24;
      17'd28160: data = 8'h22;
      17'd28161: data = 8'h1c;
      17'd28162: data = 8'h22;
      17'd28163: data = 8'h1a;
      17'd28164: data = 8'h09;
      17'd28165: data = 8'h02;
      17'd28166: data = 8'h00;
      17'd28167: data = 8'hfd;
      17'd28168: data = 8'hfc;
      17'd28169: data = 8'hf6;
      17'd28170: data = 8'hfa;
      17'd28171: data = 8'hfa;
      17'd28172: data = 8'h00;
      17'd28173: data = 8'h01;
      17'd28174: data = 8'hf4;
      17'd28175: data = 8'hfe;
      17'd28176: data = 8'hfa;
      17'd28177: data = 8'he4;
      17'd28178: data = 8'heb;
      17'd28179: data = 8'hf5;
      17'd28180: data = 8'hec;
      17'd28181: data = 8'hde;
      17'd28182: data = 8'he5;
      17'd28183: data = 8'hf5;
      17'd28184: data = 8'hf4;
      17'd28185: data = 8'hec;
      17'd28186: data = 8'hfc;
      17'd28187: data = 8'h0c;
      17'd28188: data = 8'h00;
      17'd28189: data = 8'hfd;
      17'd28190: data = 8'h06;
      17'd28191: data = 8'h0e;
      17'd28192: data = 8'hfe;
      17'd28193: data = 8'hf2;
      17'd28194: data = 8'hfc;
      17'd28195: data = 8'h04;
      17'd28196: data = 8'h01;
      17'd28197: data = 8'h00;
      17'd28198: data = 8'h0d;
      17'd28199: data = 8'h12;
      17'd28200: data = 8'h0d;
      17'd28201: data = 8'h11;
      17'd28202: data = 8'h16;
      17'd28203: data = 8'h1b;
      17'd28204: data = 8'h1c;
      17'd28205: data = 8'h15;
      17'd28206: data = 8'h1a;
      17'd28207: data = 8'h1c;
      17'd28208: data = 8'h0a;
      17'd28209: data = 8'hf9;
      17'd28210: data = 8'hf9;
      17'd28211: data = 8'h09;
      17'd28212: data = 8'h0c;
      17'd28213: data = 8'h05;
      17'd28214: data = 8'h11;
      17'd28215: data = 8'h19;
      17'd28216: data = 8'h19;
      17'd28217: data = 8'h1a;
      17'd28218: data = 8'h1a;
      17'd28219: data = 8'h11;
      17'd28220: data = 8'h09;
      17'd28221: data = 8'h05;
      17'd28222: data = 8'h0a;
      17'd28223: data = 8'h0c;
      17'd28224: data = 8'h04;
      17'd28225: data = 8'hfd;
      17'd28226: data = 8'hf9;
      17'd28227: data = 8'hfa;
      17'd28228: data = 8'hfc;
      17'd28229: data = 8'hfe;
      17'd28230: data = 8'h02;
      17'd28231: data = 8'h11;
      17'd28232: data = 8'h1b;
      17'd28233: data = 8'h1b;
      17'd28234: data = 8'h11;
      17'd28235: data = 8'h12;
      17'd28236: data = 8'h12;
      17'd28237: data = 8'h05;
      17'd28238: data = 8'hfe;
      17'd28239: data = 8'h00;
      17'd28240: data = 8'h04;
      17'd28241: data = 8'h02;
      17'd28242: data = 8'h01;
      17'd28243: data = 8'h00;
      17'd28244: data = 8'h00;
      17'd28245: data = 8'h02;
      17'd28246: data = 8'h05;
      17'd28247: data = 8'h05;
      17'd28248: data = 8'h05;
      17'd28249: data = 8'h0a;
      17'd28250: data = 8'h0c;
      17'd28251: data = 8'h0c;
      17'd28252: data = 8'h09;
      17'd28253: data = 8'h02;
      17'd28254: data = 8'hfe;
      17'd28255: data = 8'hfc;
      17'd28256: data = 8'hfa;
      17'd28257: data = 8'hfa;
      17'd28258: data = 8'hfc;
      17'd28259: data = 8'hfd;
      17'd28260: data = 8'h02;
      17'd28261: data = 8'h04;
      17'd28262: data = 8'h04;
      17'd28263: data = 8'h04;
      17'd28264: data = 8'h04;
      17'd28265: data = 8'h06;
      17'd28266: data = 8'h05;
      17'd28267: data = 8'h05;
      17'd28268: data = 8'h05;
      17'd28269: data = 8'h06;
      17'd28270: data = 8'h06;
      17'd28271: data = 8'h05;
      17'd28272: data = 8'h02;
      17'd28273: data = 8'h01;
      17'd28274: data = 8'h01;
      17'd28275: data = 8'h02;
      17'd28276: data = 8'h04;
      17'd28277: data = 8'h09;
      17'd28278: data = 8'h06;
      17'd28279: data = 8'h06;
      17'd28280: data = 8'h05;
      17'd28281: data = 8'h06;
      17'd28282: data = 8'h09;
      17'd28283: data = 8'h05;
      17'd28284: data = 8'h06;
      17'd28285: data = 8'h05;
      17'd28286: data = 8'h02;
      17'd28287: data = 8'h02;
      17'd28288: data = 8'h02;
      17'd28289: data = 8'h01;
      17'd28290: data = 8'h01;
      17'd28291: data = 8'h01;
      17'd28292: data = 8'h00;
      17'd28293: data = 8'h01;
      17'd28294: data = 8'h00;
      17'd28295: data = 8'h00;
      17'd28296: data = 8'h00;
      17'd28297: data = 8'hfe;
      17'd28298: data = 8'h00;
      17'd28299: data = 8'hfe;
      17'd28300: data = 8'hfd;
      17'd28301: data = 8'hfc;
      17'd28302: data = 8'hfa;
      17'd28303: data = 8'hfa;
      17'd28304: data = 8'hfa;
      17'd28305: data = 8'hf6;
      17'd28306: data = 8'hf5;
      17'd28307: data = 8'hf5;
      17'd28308: data = 8'hf6;
      17'd28309: data = 8'hf6;
      17'd28310: data = 8'hf6;
      17'd28311: data = 8'hf9;
      17'd28312: data = 8'hf6;
      17'd28313: data = 8'hf6;
      17'd28314: data = 8'hf5;
      17'd28315: data = 8'hf5;
      17'd28316: data = 8'hf5;
      17'd28317: data = 8'hf5;
      17'd28318: data = 8'hf5;
      17'd28319: data = 8'hf5;
      17'd28320: data = 8'hf9;
      17'd28321: data = 8'hf9;
      17'd28322: data = 8'hfa;
      17'd28323: data = 8'hf9;
      17'd28324: data = 8'hfa;
      17'd28325: data = 8'hfa;
      17'd28326: data = 8'hfa;
      17'd28327: data = 8'hfc;
      17'd28328: data = 8'hfa;
      17'd28329: data = 8'hfa;
      17'd28330: data = 8'hfc;
      17'd28331: data = 8'hfc;
      17'd28332: data = 8'hfc;
      17'd28333: data = 8'hfc;
      17'd28334: data = 8'hfc;
      17'd28335: data = 8'hfc;
      17'd28336: data = 8'hfa;
      17'd28337: data = 8'hfd;
      17'd28338: data = 8'hfa;
      17'd28339: data = 8'hf9;
      17'd28340: data = 8'hfa;
      17'd28341: data = 8'hfa;
      17'd28342: data = 8'hfa;
      17'd28343: data = 8'hf9;
      17'd28344: data = 8'hfa;
      17'd28345: data = 8'hf9;
      17'd28346: data = 8'hf9;
      17'd28347: data = 8'hf9;
      17'd28348: data = 8'hf6;
      17'd28349: data = 8'hf4;
      17'd28350: data = 8'hf2;
      17'd28351: data = 8'hf2;
      17'd28352: data = 8'hf1;
      17'd28353: data = 8'hf4;
      17'd28354: data = 8'hf4;
      17'd28355: data = 8'hf2;
      17'd28356: data = 8'hf1;
      17'd28357: data = 8'hf1;
      17'd28358: data = 8'hf2;
      17'd28359: data = 8'hf1;
      17'd28360: data = 8'hf2;
      17'd28361: data = 8'hf2;
      17'd28362: data = 8'hf4;
      17'd28363: data = 8'hf4;
      17'd28364: data = 8'hf4;
      17'd28365: data = 8'hf4;
      17'd28366: data = 8'hf5;
      17'd28367: data = 8'hf5;
      17'd28368: data = 8'hf5;
      17'd28369: data = 8'hf6;
      17'd28370: data = 8'hf6;
      17'd28371: data = 8'hf4;
      17'd28372: data = 8'hf4;
      17'd28373: data = 8'hfa;
      17'd28374: data = 8'hfc;
      17'd28375: data = 8'hfc;
      17'd28376: data = 8'hfe;
      17'd28377: data = 8'hfd;
      17'd28378: data = 8'hfe;
      17'd28379: data = 8'h00;
      17'd28380: data = 8'h00;
      17'd28381: data = 8'h00;
      17'd28382: data = 8'hfe;
      17'd28383: data = 8'hfe;
      17'd28384: data = 8'h00;
      17'd28385: data = 8'hfe;
      17'd28386: data = 8'hfe;
      17'd28387: data = 8'hfe;
      17'd28388: data = 8'hfd;
      17'd28389: data = 8'hfc;
      17'd28390: data = 8'hfc;
      17'd28391: data = 8'hfc;
      17'd28392: data = 8'hfd;
      17'd28393: data = 8'hfe;
      17'd28394: data = 8'hfe;
      17'd28395: data = 8'hfe;
      17'd28396: data = 8'hfd;
      17'd28397: data = 8'hfc;
      17'd28398: data = 8'hfc;
      17'd28399: data = 8'hfc;
      17'd28400: data = 8'hfa;
      17'd28401: data = 8'hf6;
      17'd28402: data = 8'hf6;
      17'd28403: data = 8'hfa;
      17'd28404: data = 8'hfd;
      17'd28405: data = 8'hfc;
      17'd28406: data = 8'hfc;
      17'd28407: data = 8'hfc;
      17'd28408: data = 8'hfc;
      17'd28409: data = 8'hfd;
      17'd28410: data = 8'hfe;
      17'd28411: data = 8'h00;
      17'd28412: data = 8'h00;
      17'd28413: data = 8'h00;
      17'd28414: data = 8'hfe;
      17'd28415: data = 8'hfd;
      17'd28416: data = 8'hfd;
      17'd28417: data = 8'hfc;
      17'd28418: data = 8'hfd;
      17'd28419: data = 8'h00;
      17'd28420: data = 8'h00;
      17'd28421: data = 8'h01;
      17'd28422: data = 8'h02;
      17'd28423: data = 8'h02;
      17'd28424: data = 8'h04;
      17'd28425: data = 8'h05;
      17'd28426: data = 8'h04;
      17'd28427: data = 8'h04;
      17'd28428: data = 8'h04;
      17'd28429: data = 8'h01;
      17'd28430: data = 8'h00;
      17'd28431: data = 8'h00;
      17'd28432: data = 8'h00;
      17'd28433: data = 8'h00;
      17'd28434: data = 8'h00;
      17'd28435: data = 8'h01;
      17'd28436: data = 8'h04;
      17'd28437: data = 8'h02;
      17'd28438: data = 8'h04;
      17'd28439: data = 8'h05;
      17'd28440: data = 8'h06;
      17'd28441: data = 8'h06;
      17'd28442: data = 8'h0a;
      17'd28443: data = 8'h09;
      17'd28444: data = 8'h05;
      17'd28445: data = 8'h04;
      17'd28446: data = 8'h05;
      17'd28447: data = 8'h04;
      17'd28448: data = 8'h02;
      17'd28449: data = 8'h02;
      17'd28450: data = 8'h04;
      17'd28451: data = 8'h05;
      17'd28452: data = 8'h06;
      17'd28453: data = 8'h06;
      17'd28454: data = 8'h06;
      17'd28455: data = 8'h0a;
      17'd28456: data = 8'h0a;
      17'd28457: data = 8'h0c;
      17'd28458: data = 8'h0a;
      17'd28459: data = 8'h0d;
      17'd28460: data = 8'h0d;
      17'd28461: data = 8'h0c;
      17'd28462: data = 8'h0c;
      17'd28463: data = 8'h0a;
      17'd28464: data = 8'h0c;
      17'd28465: data = 8'h0c;
      17'd28466: data = 8'h0a;
      17'd28467: data = 8'h0d;
      17'd28468: data = 8'h0e;
      17'd28469: data = 8'h11;
      17'd28470: data = 8'h13;
      17'd28471: data = 8'h15;
      17'd28472: data = 8'h16;
      17'd28473: data = 8'h16;
      17'd28474: data = 8'h16;
      17'd28475: data = 8'h15;
      17'd28476: data = 8'h15;
      17'd28477: data = 8'h15;
      17'd28478: data = 8'h15;
      17'd28479: data = 8'h11;
      17'd28480: data = 8'h12;
      17'd28481: data = 8'h12;
      17'd28482: data = 8'h11;
      17'd28483: data = 8'h0e;
      17'd28484: data = 8'h0d;
      17'd28485: data = 8'h0d;
      17'd28486: data = 8'h11;
      17'd28487: data = 8'h0d;
      17'd28488: data = 8'h0d;
      17'd28489: data = 8'h0d;
      17'd28490: data = 8'h06;
      17'd28491: data = 8'h06;
      17'd28492: data = 8'h05;
      17'd28493: data = 8'h02;
      17'd28494: data = 8'hfe;
      17'd28495: data = 8'hfe;
      17'd28496: data = 8'hfe;
      17'd28497: data = 8'hfe;
      17'd28498: data = 8'hfe;
      17'd28499: data = 8'hfd;
      17'd28500: data = 8'hfe;
      17'd28501: data = 8'hfc;
      17'd28502: data = 8'hfe;
      17'd28503: data = 8'hfd;
      17'd28504: data = 8'hfc;
      17'd28505: data = 8'hfc;
      17'd28506: data = 8'hfc;
      17'd28507: data = 8'hfc;
      17'd28508: data = 8'hfe;
      17'd28509: data = 8'hfe;
      17'd28510: data = 8'hf9;
      17'd28511: data = 8'hfa;
      17'd28512: data = 8'hfc;
      17'd28513: data = 8'hfe;
      17'd28514: data = 8'hfd;
      17'd28515: data = 8'hfe;
      17'd28516: data = 8'h01;
      17'd28517: data = 8'h02;
      17'd28518: data = 8'h06;
      17'd28519: data = 8'h05;
      17'd28520: data = 8'h05;
      17'd28521: data = 8'h04;
      17'd28522: data = 8'h04;
      17'd28523: data = 8'h04;
      17'd28524: data = 8'h05;
      17'd28525: data = 8'h04;
      17'd28526: data = 8'h04;
      17'd28527: data = 8'h04;
      17'd28528: data = 8'h04;
      17'd28529: data = 8'h04;
      17'd28530: data = 8'h04;
      17'd28531: data = 8'h02;
      17'd28532: data = 8'h04;
      17'd28533: data = 8'h06;
      17'd28534: data = 8'h05;
      17'd28535: data = 8'h04;
      17'd28536: data = 8'h04;
      17'd28537: data = 8'h00;
      17'd28538: data = 8'hfe;
      17'd28539: data = 8'hfc;
      17'd28540: data = 8'hf9;
      17'd28541: data = 8'hf6;
      17'd28542: data = 8'hf5;
      17'd28543: data = 8'hf5;
      17'd28544: data = 8'hf2;
      17'd28545: data = 8'hf1;
      17'd28546: data = 8'hf5;
      17'd28547: data = 8'hf5;
      17'd28548: data = 8'hf5;
      17'd28549: data = 8'hf4;
      17'd28550: data = 8'hf5;
      17'd28551: data = 8'hf5;
      17'd28552: data = 8'hf2;
      17'd28553: data = 8'hef;
      17'd28554: data = 8'hed;
      17'd28555: data = 8'hed;
      17'd28556: data = 8'hed;
      17'd28557: data = 8'hed;
      17'd28558: data = 8'hed;
      17'd28559: data = 8'hed;
      17'd28560: data = 8'hef;
      17'd28561: data = 8'hf2;
      17'd28562: data = 8'hf4;
      17'd28563: data = 8'hf4;
      17'd28564: data = 8'hf5;
      17'd28565: data = 8'hf5;
      17'd28566: data = 8'hf5;
      17'd28567: data = 8'hf9;
      17'd28568: data = 8'hf6;
      17'd28569: data = 8'hfc;
      17'd28570: data = 8'hf6;
      17'd28571: data = 8'hf6;
      17'd28572: data = 8'hfa;
      17'd28573: data = 8'hf9;
      17'd28574: data = 8'hfd;
      17'd28575: data = 8'hfc;
      17'd28576: data = 8'hfd;
      17'd28577: data = 8'hfe;
      17'd28578: data = 8'h00;
      17'd28579: data = 8'hfe;
      17'd28580: data = 8'h01;
      17'd28581: data = 8'h00;
      17'd28582: data = 8'hfe;
      17'd28583: data = 8'hfe;
      17'd28584: data = 8'hfe;
      17'd28585: data = 8'hfd;
      17'd28586: data = 8'hfd;
      17'd28587: data = 8'hfd;
      17'd28588: data = 8'hfd;
      17'd28589: data = 8'hfa;
      17'd28590: data = 8'hfc;
      17'd28591: data = 8'hfd;
      17'd28592: data = 8'hfc;
      17'd28593: data = 8'hfd;
      17'd28594: data = 8'hfc;
      17'd28595: data = 8'hfc;
      17'd28596: data = 8'hfc;
      17'd28597: data = 8'hfa;
      17'd28598: data = 8'hf9;
      17'd28599: data = 8'hf9;
      17'd28600: data = 8'hf6;
      17'd28601: data = 8'hf9;
      17'd28602: data = 8'hf6;
      17'd28603: data = 8'hf6;
      17'd28604: data = 8'hf5;
      17'd28605: data = 8'hf4;
      17'd28606: data = 8'hf4;
      17'd28607: data = 8'hf6;
      17'd28608: data = 8'hf6;
      17'd28609: data = 8'hf9;
      17'd28610: data = 8'hfc;
      17'd28611: data = 8'hfc;
      17'd28612: data = 8'hfe;
      17'd28613: data = 8'hfd;
      17'd28614: data = 8'hfc;
      17'd28615: data = 8'hfc;
      17'd28616: data = 8'hfa;
      17'd28617: data = 8'hfe;
      17'd28618: data = 8'hfe;
      17'd28619: data = 8'hfe;
      17'd28620: data = 8'h01;
      17'd28621: data = 8'h01;
      17'd28622: data = 8'h02;
      17'd28623: data = 8'h02;
      17'd28624: data = 8'h00;
      17'd28625: data = 8'h02;
      17'd28626: data = 8'h05;
      17'd28627: data = 8'h02;
      17'd28628: data = 8'h02;
      17'd28629: data = 8'h01;
      17'd28630: data = 8'h02;
      17'd28631: data = 8'h02;
      17'd28632: data = 8'h02;
      17'd28633: data = 8'h02;
      17'd28634: data = 8'h02;
      17'd28635: data = 8'h01;
      17'd28636: data = 8'h02;
      17'd28637: data = 8'h05;
      17'd28638: data = 8'h02;
      17'd28639: data = 8'h00;
      17'd28640: data = 8'h00;
      17'd28641: data = 8'h00;
      17'd28642: data = 8'hfe;
      17'd28643: data = 8'hfe;
      17'd28644: data = 8'hfd;
      17'd28645: data = 8'hfd;
      17'd28646: data = 8'hfd;
      17'd28647: data = 8'hfc;
      17'd28648: data = 8'h00;
      17'd28649: data = 8'hfe;
      17'd28650: data = 8'hfd;
      17'd28651: data = 8'h01;
      17'd28652: data = 8'hfe;
      17'd28653: data = 8'hfe;
      17'd28654: data = 8'hfc;
      17'd28655: data = 8'hfc;
      17'd28656: data = 8'hfc;
      17'd28657: data = 8'hf9;
      17'd28658: data = 8'hf9;
      17'd28659: data = 8'hf5;
      17'd28660: data = 8'h06;
      17'd28661: data = 8'hfe;
      17'd28662: data = 8'hfc;
      17'd28663: data = 8'h01;
      17'd28664: data = 8'hfd;
      17'd28665: data = 8'h02;
      17'd28666: data = 8'h02;
      17'd28667: data = 8'h01;
      17'd28668: data = 8'hfa;
      17'd28669: data = 8'hf9;
      17'd28670: data = 8'hfa;
      17'd28671: data = 8'hfe;
      17'd28672: data = 8'hfc;
      17'd28673: data = 8'hf9;
      17'd28674: data = 8'hfe;
      17'd28675: data = 8'h01;
      17'd28676: data = 8'h02;
      17'd28677: data = 8'h02;
      17'd28678: data = 8'hfe;
      17'd28679: data = 8'hfd;
      17'd28680: data = 8'h02;
      17'd28681: data = 8'h04;
      17'd28682: data = 8'h01;
      17'd28683: data = 8'h00;
      17'd28684: data = 8'hfd;
      17'd28685: data = 8'hfd;
      17'd28686: data = 8'hfe;
      17'd28687: data = 8'hfd;
      17'd28688: data = 8'hfc;
      17'd28689: data = 8'h00;
      17'd28690: data = 8'h00;
      17'd28691: data = 8'hfe;
      17'd28692: data = 8'h01;
      17'd28693: data = 8'h01;
      17'd28694: data = 8'h01;
      17'd28695: data = 8'h02;
      17'd28696: data = 8'h02;
      17'd28697: data = 8'h04;
      17'd28698: data = 8'h02;
      17'd28699: data = 8'h01;
      17'd28700: data = 8'h01;
      17'd28701: data = 8'h01;
      17'd28702: data = 8'hfe;
      17'd28703: data = 8'h00;
      17'd28704: data = 8'h02;
      17'd28705: data = 8'h04;
      17'd28706: data = 8'h04;
      17'd28707: data = 8'h04;
      17'd28708: data = 8'h06;
      17'd28709: data = 8'h0a;
      17'd28710: data = 8'h0a;
      17'd28711: data = 8'h09;
      17'd28712: data = 8'h09;
      17'd28713: data = 8'h06;
      17'd28714: data = 8'h06;
      17'd28715: data = 8'h06;
      17'd28716: data = 8'h05;
      17'd28717: data = 8'h06;
      17'd28718: data = 8'h09;
      17'd28719: data = 8'h09;
      17'd28720: data = 8'h06;
      17'd28721: data = 8'h09;
      17'd28722: data = 8'h05;
      17'd28723: data = 8'h06;
      17'd28724: data = 8'h06;
      17'd28725: data = 8'h05;
      17'd28726: data = 8'h09;
      17'd28727: data = 8'h06;
      17'd28728: data = 8'h05;
      17'd28729: data = 8'h06;
      17'd28730: data = 8'h04;
      17'd28731: data = 8'h04;
      17'd28732: data = 8'h05;
      17'd28733: data = 8'h01;
      17'd28734: data = 8'h01;
      17'd28735: data = 8'h04;
      17'd28736: data = 8'h02;
      17'd28737: data = 8'h01;
      17'd28738: data = 8'h02;
      17'd28739: data = 8'h02;
      17'd28740: data = 8'h02;
      17'd28741: data = 8'h01;
      17'd28742: data = 8'h01;
      17'd28743: data = 8'h01;
      17'd28744: data = 8'h01;
      17'd28745: data = 8'h02;
      17'd28746: data = 8'h02;
      17'd28747: data = 8'h01;
      17'd28748: data = 8'h01;
      17'd28749: data = 8'h01;
      17'd28750: data = 8'h00;
      17'd28751: data = 8'h00;
      17'd28752: data = 8'h01;
      17'd28753: data = 8'h04;
      17'd28754: data = 8'h04;
      17'd28755: data = 8'h05;
      17'd28756: data = 8'h09;
      17'd28757: data = 8'h06;
      17'd28758: data = 8'h09;
      17'd28759: data = 8'h09;
      17'd28760: data = 8'h09;
      17'd28761: data = 8'h06;
      17'd28762: data = 8'h06;
      17'd28763: data = 8'h05;
      17'd28764: data = 8'h04;
      17'd28765: data = 8'h05;
      17'd28766: data = 8'h04;
      17'd28767: data = 8'h02;
      17'd28768: data = 8'h04;
      17'd28769: data = 8'h05;
      17'd28770: data = 8'h02;
      17'd28771: data = 8'h02;
      17'd28772: data = 8'h02;
      17'd28773: data = 8'h04;
      17'd28774: data = 8'h01;
      17'd28775: data = 8'h01;
      17'd28776: data = 8'h00;
      17'd28777: data = 8'hfd;
      17'd28778: data = 8'hfa;
      17'd28779: data = 8'hf9;
      17'd28780: data = 8'hfd;
      17'd28781: data = 8'hfd;
      17'd28782: data = 8'hfc;
      17'd28783: data = 8'hfe;
      17'd28784: data = 8'h00;
      17'd28785: data = 8'hfd;
      17'd28786: data = 8'hfd;
      17'd28787: data = 8'hfd;
      17'd28788: data = 8'hfa;
      17'd28789: data = 8'hf9;
      17'd28790: data = 8'hfc;
      17'd28791: data = 8'hf9;
      17'd28792: data = 8'hf6;
      17'd28793: data = 8'hf6;
      17'd28794: data = 8'hf9;
      17'd28795: data = 8'hf9;
      17'd28796: data = 8'hf5;
      17'd28797: data = 8'hf6;
      17'd28798: data = 8'hf9;
      17'd28799: data = 8'hf9;
      17'd28800: data = 8'hfa;
      17'd28801: data = 8'hfa;
      17'd28802: data = 8'hf9;
      17'd28803: data = 8'hfc;
      17'd28804: data = 8'hfc;
      17'd28805: data = 8'hfa;
      17'd28806: data = 8'hfd;
      17'd28807: data = 8'hfc;
      17'd28808: data = 8'hfd;
      17'd28809: data = 8'hfa;
      17'd28810: data = 8'hf6;
      17'd28811: data = 8'hfa;
      17'd28812: data = 8'hf9;
      17'd28813: data = 8'hf9;
      17'd28814: data = 8'hfa;
      17'd28815: data = 8'hfa;
      17'd28816: data = 8'hfc;
      17'd28817: data = 8'hfd;
      17'd28818: data = 8'hfe;
      17'd28819: data = 8'h00;
      17'd28820: data = 8'h00;
      17'd28821: data = 8'hfe;
      17'd28822: data = 8'hfc;
      17'd28823: data = 8'hfc;
      17'd28824: data = 8'hfa;
      17'd28825: data = 8'hf9;
      17'd28826: data = 8'hfa;
      17'd28827: data = 8'hfc;
      17'd28828: data = 8'hfc;
      17'd28829: data = 8'hfd;
      17'd28830: data = 8'hfd;
      17'd28831: data = 8'hfc;
      17'd28832: data = 8'hfc;
      17'd28833: data = 8'hfe;
      17'd28834: data = 8'hfd;
      17'd28835: data = 8'hfd;
      17'd28836: data = 8'hfe;
      17'd28837: data = 8'hfd;
      17'd28838: data = 8'hfe;
      17'd28839: data = 8'hfd;
      17'd28840: data = 8'hfd;
      17'd28841: data = 8'hfc;
      17'd28842: data = 8'hfc;
      17'd28843: data = 8'hfa;
      17'd28844: data = 8'hf9;
      17'd28845: data = 8'hf9;
      17'd28846: data = 8'hf9;
      17'd28847: data = 8'hf6;
      17'd28848: data = 8'hf9;
      17'd28849: data = 8'hf6;
      17'd28850: data = 8'hf6;
      17'd28851: data = 8'hf6;
      17'd28852: data = 8'hfa;
      17'd28853: data = 8'hf5;
      17'd28854: data = 8'hf5;
      17'd28855: data = 8'hf9;
      17'd28856: data = 8'hf5;
      17'd28857: data = 8'hf6;
      17'd28858: data = 8'hf5;
      17'd28859: data = 8'hf4;
      17'd28860: data = 8'hf5;
      17'd28861: data = 8'hf5;
      17'd28862: data = 8'hf2;
      17'd28863: data = 8'hf2;
      17'd28864: data = 8'hf2;
      17'd28865: data = 8'hf4;
      17'd28866: data = 8'hf5;
      17'd28867: data = 8'hf9;
      17'd28868: data = 8'hfc;
      17'd28869: data = 8'hfc;
      17'd28870: data = 8'hfe;
      17'd28871: data = 8'hfe;
      17'd28872: data = 8'h00;
      17'd28873: data = 8'h01;
      17'd28874: data = 8'hfe;
      17'd28875: data = 8'hfe;
      17'd28876: data = 8'hfe;
      17'd28877: data = 8'hfc;
      17'd28878: data = 8'hf9;
      17'd28879: data = 8'hfa;
      17'd28880: data = 8'hf9;
      17'd28881: data = 8'hf9;
      17'd28882: data = 8'hfa;
      17'd28883: data = 8'hfd;
      17'd28884: data = 8'hfe;
      17'd28885: data = 8'hfd;
      17'd28886: data = 8'h00;
      17'd28887: data = 8'hfe;
      17'd28888: data = 8'hfd;
      17'd28889: data = 8'hfd;
      17'd28890: data = 8'hfa;
      17'd28891: data = 8'hf9;
      17'd28892: data = 8'hf9;
      17'd28893: data = 8'hf9;
      17'd28894: data = 8'hf9;
      17'd28895: data = 8'hfa;
      17'd28896: data = 8'hfa;
      17'd28897: data = 8'hf9;
      17'd28898: data = 8'hfd;
      17'd28899: data = 8'hfd;
      17'd28900: data = 8'hfd;
      17'd28901: data = 8'hfd;
      17'd28902: data = 8'hfa;
      17'd28903: data = 8'hf9;
      17'd28904: data = 8'hf9;
      17'd28905: data = 8'hf6;
      17'd28906: data = 8'hf4;
      17'd28907: data = 8'hf1;
      17'd28908: data = 8'hef;
      17'd28909: data = 8'hf2;
      17'd28910: data = 8'hf2;
      17'd28911: data = 8'hf2;
      17'd28912: data = 8'hf6;
      17'd28913: data = 8'hfa;
      17'd28914: data = 8'hfc;
      17'd28915: data = 8'hfc;
      17'd28916: data = 8'hfc;
      17'd28917: data = 8'hfd;
      17'd28918: data = 8'hfe;
      17'd28919: data = 8'hfe;
      17'd28920: data = 8'hfe;
      17'd28921: data = 8'h01;
      17'd28922: data = 8'h00;
      17'd28923: data = 8'hfe;
      17'd28924: data = 8'h00;
      17'd28925: data = 8'h00;
      17'd28926: data = 8'h01;
      17'd28927: data = 8'h01;
      17'd28928: data = 8'h04;
      17'd28929: data = 8'h06;
      17'd28930: data = 8'h06;
      17'd28931: data = 8'h0a;
      17'd28932: data = 8'h0a;
      17'd28933: data = 8'h09;
      17'd28934: data = 8'h0a;
      17'd28935: data = 8'h09;
      17'd28936: data = 8'h09;
      17'd28937: data = 8'h06;
      17'd28938: data = 8'h05;
      17'd28939: data = 8'h06;
      17'd28940: data = 8'h05;
      17'd28941: data = 8'h06;
      17'd28942: data = 8'h06;
      17'd28943: data = 8'h05;
      17'd28944: data = 8'h05;
      17'd28945: data = 8'h09;
      17'd28946: data = 8'h09;
      17'd28947: data = 8'h09;
      17'd28948: data = 8'h09;
      17'd28949: data = 8'h09;
      17'd28950: data = 8'h06;
      17'd28951: data = 8'h06;
      17'd28952: data = 8'h06;
      17'd28953: data = 8'h04;
      17'd28954: data = 8'h01;
      17'd28955: data = 8'h01;
      17'd28956: data = 8'h02;
      17'd28957: data = 8'h02;
      17'd28958: data = 8'h01;
      17'd28959: data = 8'h02;
      17'd28960: data = 8'h02;
      17'd28961: data = 8'h04;
      17'd28962: data = 8'h04;
      17'd28963: data = 8'h05;
      17'd28964: data = 8'h05;
      17'd28965: data = 8'h02;
      17'd28966: data = 8'h02;
      17'd28967: data = 8'h01;
      17'd28968: data = 8'h02;
      17'd28969: data = 8'h00;
      17'd28970: data = 8'hfe;
      17'd28971: data = 8'h01;
      17'd28972: data = 8'h02;
      17'd28973: data = 8'h01;
      17'd28974: data = 8'h02;
      17'd28975: data = 8'h05;
      17'd28976: data = 8'h06;
      17'd28977: data = 8'h09;
      17'd28978: data = 8'h06;
      17'd28979: data = 8'h06;
      17'd28980: data = 8'h06;
      17'd28981: data = 8'h05;
      17'd28982: data = 8'h06;
      17'd28983: data = 8'h09;
      17'd28984: data = 8'h06;
      17'd28985: data = 8'h09;
      17'd28986: data = 8'h05;
      17'd28987: data = 8'h06;
      17'd28988: data = 8'h09;
      17'd28989: data = 8'h0a;
      17'd28990: data = 8'h0c;
      17'd28991: data = 8'h0c;
      17'd28992: data = 8'h0d;
      17'd28993: data = 8'h0e;
      17'd28994: data = 8'h0a;
      17'd28995: data = 8'h09;
      17'd28996: data = 8'h06;
      17'd28997: data = 8'h06;
      17'd28998: data = 8'h05;
      17'd28999: data = 8'h04;
      17'd29000: data = 8'h04;
      17'd29001: data = 8'h02;
      17'd29002: data = 8'h02;
      17'd29003: data = 8'h01;
      17'd29004: data = 8'h00;
      17'd29005: data = 8'h00;
      17'd29006: data = 8'h01;
      17'd29007: data = 8'h00;
      17'd29008: data = 8'h00;
      17'd29009: data = 8'h00;
      17'd29010: data = 8'hfe;
      17'd29011: data = 8'hfe;
      17'd29012: data = 8'hfd;
      17'd29013: data = 8'hfc;
      17'd29014: data = 8'hfa;
      17'd29015: data = 8'hfa;
      17'd29016: data = 8'hf9;
      17'd29017: data = 8'hf6;
      17'd29018: data = 8'hf6;
      17'd29019: data = 8'hf6;
      17'd29020: data = 8'hfa;
      17'd29021: data = 8'hfc;
      17'd29022: data = 8'hfc;
      17'd29023: data = 8'hfe;
      17'd29024: data = 8'hfd;
      17'd29025: data = 8'hfd;
      17'd29026: data = 8'h00;
      17'd29027: data = 8'hfe;
      17'd29028: data = 8'h00;
      17'd29029: data = 8'h01;
      17'd29030: data = 8'h02;
      17'd29031: data = 8'h02;
      17'd29032: data = 8'h02;
      17'd29033: data = 8'h02;
      17'd29034: data = 8'h02;
      17'd29035: data = 8'h02;
      17'd29036: data = 8'h04;
      17'd29037: data = 8'h05;
      17'd29038: data = 8'h05;
      17'd29039: data = 8'h05;
      17'd29040: data = 8'h05;
      17'd29041: data = 8'h04;
      17'd29042: data = 8'h04;
      17'd29043: data = 8'h02;
      17'd29044: data = 8'h01;
      17'd29045: data = 8'h00;
      17'd29046: data = 8'hfd;
      17'd29047: data = 8'hfd;
      17'd29048: data = 8'hfd;
      17'd29049: data = 8'hfc;
      17'd29050: data = 8'hfc;
      17'd29051: data = 8'hfc;
      17'd29052: data = 8'hfa;
      17'd29053: data = 8'hfc;
      17'd29054: data = 8'hfe;
      17'd29055: data = 8'hfd;
      17'd29056: data = 8'hfd;
      17'd29057: data = 8'hfe;
      17'd29058: data = 8'hfc;
      17'd29059: data = 8'hfa;
      17'd29060: data = 8'hf9;
      17'd29061: data = 8'hf6;
      17'd29062: data = 8'hf5;
      17'd29063: data = 8'hf4;
      17'd29064: data = 8'hf5;
      17'd29065: data = 8'hf9;
      17'd29066: data = 8'hf9;
      17'd29067: data = 8'hfa;
      17'd29068: data = 8'hfa;
      17'd29069: data = 8'hfc;
      17'd29070: data = 8'hfc;
      17'd29071: data = 8'hfa;
      17'd29072: data = 8'hfc;
      17'd29073: data = 8'hfc;
      17'd29074: data = 8'hfc;
      17'd29075: data = 8'hfc;
      17'd29076: data = 8'hfc;
      17'd29077: data = 8'hfc;
      17'd29078: data = 8'hfc;
      17'd29079: data = 8'hfd;
      17'd29080: data = 8'hfc;
      17'd29081: data = 8'hfd;
      17'd29082: data = 8'hfe;
      17'd29083: data = 8'h00;
      17'd29084: data = 8'h02;
      17'd29085: data = 8'h01;
      17'd29086: data = 8'h01;
      17'd29087: data = 8'h00;
      17'd29088: data = 8'h00;
      17'd29089: data = 8'hfd;
      17'd29090: data = 8'hfd;
      17'd29091: data = 8'hfd;
      17'd29092: data = 8'hfa;
      17'd29093: data = 8'hfc;
      17'd29094: data = 8'hfc;
      17'd29095: data = 8'hfa;
      17'd29096: data = 8'hfc;
      17'd29097: data = 8'hfd;
      17'd29098: data = 8'hfc;
      17'd29099: data = 8'hfa;
      17'd29100: data = 8'hfc;
      17'd29101: data = 8'hfc;
      17'd29102: data = 8'hfc;
      17'd29103: data = 8'hfc;
      17'd29104: data = 8'hfc;
      17'd29105: data = 8'hfc;
      17'd29106: data = 8'hfc;
      17'd29107: data = 8'hfa;
      17'd29108: data = 8'hfa;
      17'd29109: data = 8'hf9;
      17'd29110: data = 8'hf9;
      17'd29111: data = 8'hf9;
      17'd29112: data = 8'hfa;
      17'd29113: data = 8'hf9;
      17'd29114: data = 8'hfa;
      17'd29115: data = 8'hfa;
      17'd29116: data = 8'hf9;
      17'd29117: data = 8'hfa;
      17'd29118: data = 8'hfc;
      17'd29119: data = 8'hfc;
      17'd29120: data = 8'hfc;
      17'd29121: data = 8'hfd;
      17'd29122: data = 8'hfe;
      17'd29123: data = 8'hfe;
      17'd29124: data = 8'h00;
      17'd29125: data = 8'h00;
      17'd29126: data = 8'hfe;
      17'd29127: data = 8'hfd;
      17'd29128: data = 8'hfd;
      17'd29129: data = 8'hfd;
      17'd29130: data = 8'hfd;
      17'd29131: data = 8'hfc;
      17'd29132: data = 8'hfa;
      17'd29133: data = 8'hfc;
      17'd29134: data = 8'hfd;
      17'd29135: data = 8'hfc;
      17'd29136: data = 8'hfc;
      17'd29137: data = 8'hfd;
      17'd29138: data = 8'hfe;
      17'd29139: data = 8'hfd;
      17'd29140: data = 8'hfd;
      17'd29141: data = 8'hfd;
      17'd29142: data = 8'hfa;
      17'd29143: data = 8'hf9;
      17'd29144: data = 8'hf6;
      17'd29145: data = 8'hf9;
      17'd29146: data = 8'hfa;
      17'd29147: data = 8'hfa;
      17'd29148: data = 8'hfa;
      17'd29149: data = 8'hfc;
      17'd29150: data = 8'hfc;
      17'd29151: data = 8'hfd;
      17'd29152: data = 8'h00;
      17'd29153: data = 8'h00;
      17'd29154: data = 8'h01;
      17'd29155: data = 8'h01;
      17'd29156: data = 8'h00;
      17'd29157: data = 8'h01;
      17'd29158: data = 8'h01;
      17'd29159: data = 8'h00;
      17'd29160: data = 8'h00;
      17'd29161: data = 8'hfe;
      17'd29162: data = 8'h00;
      17'd29163: data = 8'h00;
      17'd29164: data = 8'h00;
      17'd29165: data = 8'h02;
      17'd29166: data = 8'h04;
      17'd29167: data = 8'h05;
      17'd29168: data = 8'h05;
      17'd29169: data = 8'h06;
      17'd29170: data = 8'h06;
      17'd29171: data = 8'h05;
      17'd29172: data = 8'h05;
      17'd29173: data = 8'h05;
      17'd29174: data = 8'h05;
      17'd29175: data = 8'h02;
      17'd29176: data = 8'h04;
      17'd29177: data = 8'h04;
      17'd29178: data = 8'h02;
      17'd29179: data = 8'h04;
      17'd29180: data = 8'h02;
      17'd29181: data = 8'h05;
      17'd29182: data = 8'h05;
      17'd29183: data = 8'h05;
      17'd29184: data = 8'h05;
      17'd29185: data = 8'h04;
      17'd29186: data = 8'h02;
      17'd29187: data = 8'h02;
      17'd29188: data = 8'h01;
      17'd29189: data = 8'h00;
      17'd29190: data = 8'h00;
      17'd29191: data = 8'h00;
      17'd29192: data = 8'h01;
      17'd29193: data = 8'h00;
      17'd29194: data = 8'h01;
      17'd29195: data = 8'h04;
      17'd29196: data = 8'h04;
      17'd29197: data = 8'h04;
      17'd29198: data = 8'h04;
      17'd29199: data = 8'h05;
      17'd29200: data = 8'h01;
      17'd29201: data = 8'h01;
      17'd29202: data = 8'h01;
      17'd29203: data = 8'h01;
      17'd29204: data = 8'h00;
      17'd29205: data = 8'hfd;
      17'd29206: data = 8'hfe;
      17'd29207: data = 8'hfe;
      17'd29208: data = 8'hfe;
      17'd29209: data = 8'h00;
      17'd29210: data = 8'h02;
      17'd29211: data = 8'h02;
      17'd29212: data = 8'h01;
      17'd29213: data = 8'h01;
      17'd29214: data = 8'h02;
      17'd29215: data = 8'h00;
      17'd29216: data = 8'h01;
      17'd29217: data = 8'h01;
      17'd29218: data = 8'h00;
      17'd29219: data = 8'h00;
      17'd29220: data = 8'h00;
      17'd29221: data = 8'h00;
      17'd29222: data = 8'h00;
      17'd29223: data = 8'h01;
      17'd29224: data = 8'h01;
      17'd29225: data = 8'h02;
      17'd29226: data = 8'h02;
      17'd29227: data = 8'h02;
      17'd29228: data = 8'h04;
      17'd29229: data = 8'h05;
      17'd29230: data = 8'h04;
      17'd29231: data = 8'h02;
      17'd29232: data = 8'h05;
      17'd29233: data = 8'h05;
      17'd29234: data = 8'h02;
      17'd29235: data = 8'h02;
      17'd29236: data = 8'h04;
      17'd29237: data = 8'h02;
      17'd29238: data = 8'h01;
      17'd29239: data = 8'h01;
      17'd29240: data = 8'h00;
      17'd29241: data = 8'h00;
      17'd29242: data = 8'h00;
      17'd29243: data = 8'h00;
      17'd29244: data = 8'h00;
      17'd29245: data = 8'h00;
      17'd29246: data = 8'h00;
      17'd29247: data = 8'hfe;
      17'd29248: data = 8'h00;
      17'd29249: data = 8'hfd;
      17'd29250: data = 8'hfc;
      17'd29251: data = 8'hfc;
      17'd29252: data = 8'hfa;
      17'd29253: data = 8'hfa;
      17'd29254: data = 8'hfc;
      17'd29255: data = 8'hfd;
      17'd29256: data = 8'hfd;
      17'd29257: data = 8'hfd;
      17'd29258: data = 8'hfc;
      17'd29259: data = 8'hfd;
      17'd29260: data = 8'hfd;
      17'd29261: data = 8'hfd;
      17'd29262: data = 8'hfe;
      17'd29263: data = 8'h00;
      17'd29264: data = 8'h01;
      17'd29265: data = 8'h00;
      17'd29266: data = 8'h01;
      17'd29267: data = 8'h01;
      17'd29268: data = 8'h01;
      17'd29269: data = 8'h02;
      17'd29270: data = 8'h01;
      17'd29271: data = 8'h02;
      17'd29272: data = 8'h01;
      17'd29273: data = 8'h02;
      17'd29274: data = 8'h04;
      17'd29275: data = 8'h04;
      17'd29276: data = 8'h05;
      17'd29277: data = 8'h04;
      17'd29278: data = 8'h04;
      17'd29279: data = 8'h01;
      17'd29280: data = 8'h01;
      17'd29281: data = 8'h01;
      17'd29282: data = 8'h00;
      17'd29283: data = 8'hfe;
      17'd29284: data = 8'h00;
      17'd29285: data = 8'h01;
      17'd29286: data = 8'h00;
      17'd29287: data = 8'h00;
      17'd29288: data = 8'h00;
      17'd29289: data = 8'h00;
      17'd29290: data = 8'h00;
      17'd29291: data = 8'h01;
      17'd29292: data = 8'h00;
      17'd29293: data = 8'hfd;
      17'd29294: data = 8'hfe;
      17'd29295: data = 8'hfc;
      17'd29296: data = 8'hfd;
      17'd29297: data = 8'hfd;
      17'd29298: data = 8'hfc;
      17'd29299: data = 8'hfc;
      17'd29300: data = 8'hfc;
      17'd29301: data = 8'hfc;
      17'd29302: data = 8'hfc;
      17'd29303: data = 8'hfc;
      17'd29304: data = 8'hfd;
      17'd29305: data = 8'hfd;
      17'd29306: data = 8'hfe;
      17'd29307: data = 8'hfe;
      17'd29308: data = 8'hfe;
      17'd29309: data = 8'hfe;
      17'd29310: data = 8'hfe;
      17'd29311: data = 8'h00;
      17'd29312: data = 8'h00;
      17'd29313: data = 8'h00;
      17'd29314: data = 8'h01;
      17'd29315: data = 8'h00;
      17'd29316: data = 8'h00;
      17'd29317: data = 8'h00;
      17'd29318: data = 8'hfe;
      17'd29319: data = 8'h00;
      17'd29320: data = 8'h01;
      17'd29321: data = 8'h01;
      17'd29322: data = 8'h01;
      17'd29323: data = 8'h00;
      17'd29324: data = 8'h01;
      17'd29325: data = 8'h01;
      17'd29326: data = 8'h00;
      17'd29327: data = 8'h00;
      17'd29328: data = 8'h01;
      17'd29329: data = 8'h00;
      17'd29330: data = 8'h00;
      17'd29331: data = 8'hfe;
      17'd29332: data = 8'hfd;
      17'd29333: data = 8'hfe;
      17'd29334: data = 8'hfe;
      17'd29335: data = 8'hfe;
      17'd29336: data = 8'hfe;
      17'd29337: data = 8'hfe;
      17'd29338: data = 8'hfe;
      17'd29339: data = 8'h00;
      17'd29340: data = 8'h00;
      17'd29341: data = 8'hfe;
      17'd29342: data = 8'h00;
      17'd29343: data = 8'h00;
      17'd29344: data = 8'h00;
      17'd29345: data = 8'hfe;
      17'd29346: data = 8'hfe;
      17'd29347: data = 8'h00;
      17'd29348: data = 8'hfe;
      17'd29349: data = 8'hfe;
      17'd29350: data = 8'hfd;
      17'd29351: data = 8'hfd;
      17'd29352: data = 8'hfe;
      17'd29353: data = 8'hfe;
      17'd29354: data = 8'h00;
      17'd29355: data = 8'h01;
      17'd29356: data = 8'h01;
      17'd29357: data = 8'h00;
      17'd29358: data = 8'h02;
      17'd29359: data = 8'h00;
      17'd29360: data = 8'hfe;
      17'd29361: data = 8'h01;
      17'd29362: data = 8'h00;
      17'd29363: data = 8'h00;
      17'd29364: data = 8'h00;
      17'd29365: data = 8'hfe;
      17'd29366: data = 8'hfe;
      17'd29367: data = 8'hfe;
      17'd29368: data = 8'hfd;
      17'd29369: data = 8'h00;
      17'd29370: data = 8'h01;
      17'd29371: data = 8'hfe;
      17'd29372: data = 8'hfe;
      17'd29373: data = 8'h00;
      17'd29374: data = 8'h00;
      17'd29375: data = 8'hfe;
      17'd29376: data = 8'h01;
      17'd29377: data = 8'h00;
      17'd29378: data = 8'hfd;
      17'd29379: data = 8'hfe;
      17'd29380: data = 8'hfe;
      17'd29381: data = 8'hfd;
      17'd29382: data = 8'hfd;
      17'd29383: data = 8'hfe;
      17'd29384: data = 8'h00;
      17'd29385: data = 8'hfe;
      17'd29386: data = 8'hfe;
      17'd29387: data = 8'h00;
      17'd29388: data = 8'h00;
      17'd29389: data = 8'h00;
      17'd29390: data = 8'h00;
      17'd29391: data = 8'h00;
      17'd29392: data = 8'h00;
      17'd29393: data = 8'h00;
      17'd29394: data = 8'h01;
      17'd29395: data = 8'h01;
      17'd29396: data = 8'h01;
      17'd29397: data = 8'h04;
      17'd29398: data = 8'h05;
      17'd29399: data = 8'h04;
      17'd29400: data = 8'h04;
      17'd29401: data = 8'h04;
      17'd29402: data = 8'h02;
      17'd29403: data = 8'h02;
      17'd29404: data = 8'h04;
      17'd29405: data = 8'h04;
      17'd29406: data = 8'h01;
      17'd29407: data = 8'h02;
      17'd29408: data = 8'h00;
      17'd29409: data = 8'h00;
      17'd29410: data = 8'h00;
      17'd29411: data = 8'h01;
      17'd29412: data = 8'h02;
      17'd29413: data = 8'h00;
      17'd29414: data = 8'h00;
      17'd29415: data = 8'h01;
      17'd29416: data = 8'h02;
      17'd29417: data = 8'h01;
      17'd29418: data = 8'h00;
      17'd29419: data = 8'h01;
      17'd29420: data = 8'h00;
      17'd29421: data = 8'hfd;
      17'd29422: data = 8'hfc;
      17'd29423: data = 8'hfc;
      17'd29424: data = 8'hfa;
      17'd29425: data = 8'hfd;
      17'd29426: data = 8'hfe;
      17'd29427: data = 8'hfe;
      17'd29428: data = 8'hfd;
      17'd29429: data = 8'h00;
      17'd29430: data = 8'h00;
      17'd29431: data = 8'h00;
      17'd29432: data = 8'h01;
      17'd29433: data = 8'h01;
      17'd29434: data = 8'h02;
      17'd29435: data = 8'h02;
      17'd29436: data = 8'h02;
      17'd29437: data = 8'h02;
      17'd29438: data = 8'h00;
      17'd29439: data = 8'h00;
      17'd29440: data = 8'h00;
      17'd29441: data = 8'h01;
      17'd29442: data = 8'h01;
      17'd29443: data = 8'h01;
      17'd29444: data = 8'h01;
      17'd29445: data = 8'h02;
      17'd29446: data = 8'h04;
      17'd29447: data = 8'h02;
      17'd29448: data = 8'h04;
      17'd29449: data = 8'h02;
      17'd29450: data = 8'h01;
      17'd29451: data = 8'h02;
      17'd29452: data = 8'h00;
      17'd29453: data = 8'hfe;
      17'd29454: data = 8'h00;
      17'd29455: data = 8'hfe;
      17'd29456: data = 8'h00;
      17'd29457: data = 8'hfe;
      17'd29458: data = 8'hfc;
      17'd29459: data = 8'hfd;
      17'd29460: data = 8'hfd;
      17'd29461: data = 8'hfd;
      17'd29462: data = 8'hfe;
      17'd29463: data = 8'hfe;
      17'd29464: data = 8'hfe;
      17'd29465: data = 8'hfd;
      17'd29466: data = 8'hfe;
      17'd29467: data = 8'hfd;
      17'd29468: data = 8'hfd;
      17'd29469: data = 8'hfd;
      17'd29470: data = 8'hfc;
      17'd29471: data = 8'hfd;
      17'd29472: data = 8'hfd;
      17'd29473: data = 8'hfd;
      17'd29474: data = 8'hfe;
      17'd29475: data = 8'hfe;
      17'd29476: data = 8'hfc;
      17'd29477: data = 8'hfd;
      17'd29478: data = 8'hfd;
      17'd29479: data = 8'hfa;
      17'd29480: data = 8'hfc;
      17'd29481: data = 8'hfd;
      17'd29482: data = 8'hfa;
      17'd29483: data = 8'hfa;
      17'd29484: data = 8'hfc;
      17'd29485: data = 8'hfd;
      17'd29486: data = 8'hfc;
      17'd29487: data = 8'hfc;
      17'd29488: data = 8'hfc;
      17'd29489: data = 8'hfc;
      17'd29490: data = 8'hfc;
      17'd29491: data = 8'hfc;
      17'd29492: data = 8'hfc;
      17'd29493: data = 8'hfc;
      17'd29494: data = 8'hfc;
      17'd29495: data = 8'hfc;
      17'd29496: data = 8'hfd;
      17'd29497: data = 8'hfc;
      17'd29498: data = 8'hfe;
      17'd29499: data = 8'h00;
      17'd29500: data = 8'h00;
      17'd29501: data = 8'h01;
      17'd29502: data = 8'h01;
      17'd29503: data = 8'h02;
      17'd29504: data = 8'h02;
      17'd29505: data = 8'h01;
      17'd29506: data = 8'h00;
      17'd29507: data = 8'h00;
      17'd29508: data = 8'h01;
      17'd29509: data = 8'h01;
      17'd29510: data = 8'hfe;
      17'd29511: data = 8'hfd;
      17'd29512: data = 8'hfd;
      17'd29513: data = 8'hfe;
      17'd29514: data = 8'h00;
      17'd29515: data = 8'h00;
      17'd29516: data = 8'h00;
      17'd29517: data = 8'hfe;
      17'd29518: data = 8'h00;
      17'd29519: data = 8'hfe;
      17'd29520: data = 8'hfd;
      17'd29521: data = 8'hfd;
      17'd29522: data = 8'hfd;
      17'd29523: data = 8'hfa;
      17'd29524: data = 8'hfd;
      17'd29525: data = 8'hfc;
      17'd29526: data = 8'hfd;
      17'd29527: data = 8'hfc;
      17'd29528: data = 8'hf9;
      17'd29529: data = 8'hf9;
      17'd29530: data = 8'hf9;
      17'd29531: data = 8'hf9;
      17'd29532: data = 8'hf9;
      17'd29533: data = 8'hfa;
      17'd29534: data = 8'hfa;
      17'd29535: data = 8'hfc;
      17'd29536: data = 8'hfc;
      17'd29537: data = 8'hfd;
      17'd29538: data = 8'hfe;
      17'd29539: data = 8'hfe;
      17'd29540: data = 8'hfe;
      17'd29541: data = 8'hfe;
      17'd29542: data = 8'hfe;
      17'd29543: data = 8'hfe;
      17'd29544: data = 8'hfe;
      17'd29545: data = 8'hfe;
      17'd29546: data = 8'hfe;
      17'd29547: data = 8'hfd;
      17'd29548: data = 8'h00;
      17'd29549: data = 8'h01;
      17'd29550: data = 8'h02;
      17'd29551: data = 8'h04;
      17'd29552: data = 8'h04;
      17'd29553: data = 8'h02;
      17'd29554: data = 8'h04;
      17'd29555: data = 8'h02;
      17'd29556: data = 8'h01;
      17'd29557: data = 8'h00;
      17'd29558: data = 8'hfe;
      17'd29559: data = 8'h01;
      17'd29560: data = 8'h01;
      17'd29561: data = 8'h01;
      17'd29562: data = 8'h02;
      17'd29563: data = 8'h02;
      17'd29564: data = 8'h02;
      17'd29565: data = 8'h02;
      17'd29566: data = 8'h01;
      17'd29567: data = 8'h00;
      17'd29568: data = 8'h00;
      17'd29569: data = 8'hfd;
      17'd29570: data = 8'hfd;
      17'd29571: data = 8'hfd;
      17'd29572: data = 8'hf9;
      17'd29573: data = 8'hfa;
      17'd29574: data = 8'hfa;
      17'd29575: data = 8'hfa;
      17'd29576: data = 8'hfd;
      17'd29577: data = 8'hfe;
      17'd29578: data = 8'hfe;
      17'd29579: data = 8'h00;
      17'd29580: data = 8'h00;
      17'd29581: data = 8'h00;
      17'd29582: data = 8'hfe;
      17'd29583: data = 8'hfe;
      17'd29584: data = 8'hfd;
      17'd29585: data = 8'hfa;
      17'd29586: data = 8'hfc;
      17'd29587: data = 8'hfc;
      17'd29588: data = 8'hfc;
      17'd29589: data = 8'hfc;
      17'd29590: data = 8'hfc;
      17'd29591: data = 8'hfd;
      17'd29592: data = 8'hfe;
      17'd29593: data = 8'h01;
      17'd29594: data = 8'h04;
      17'd29595: data = 8'h04;
      17'd29596: data = 8'h05;
      17'd29597: data = 8'h05;
      17'd29598: data = 8'h04;
      17'd29599: data = 8'h05;
      17'd29600: data = 8'h04;
      17'd29601: data = 8'h01;
      17'd29602: data = 8'h00;
      17'd29603: data = 8'h00;
      17'd29604: data = 8'h00;
      17'd29605: data = 8'h00;
      17'd29606: data = 8'h01;
      17'd29607: data = 8'h02;
      17'd29608: data = 8'h02;
      17'd29609: data = 8'h02;
      17'd29610: data = 8'h04;
      17'd29611: data = 8'h04;
      17'd29612: data = 8'h04;
      17'd29613: data = 8'h04;
      17'd29614: data = 8'h02;
      17'd29615: data = 8'h01;
      17'd29616: data = 8'h01;
      17'd29617: data = 8'hfe;
      17'd29618: data = 8'hfc;
      17'd29619: data = 8'hfa;
      17'd29620: data = 8'hf9;
      17'd29621: data = 8'hf9;
      17'd29622: data = 8'hfa;
      17'd29623: data = 8'hfc;
      17'd29624: data = 8'hfc;
      17'd29625: data = 8'hfd;
      17'd29626: data = 8'h00;
      17'd29627: data = 8'h00;
      17'd29628: data = 8'h01;
      17'd29629: data = 8'h00;
      17'd29630: data = 8'h00;
      17'd29631: data = 8'h00;
      17'd29632: data = 8'h01;
      17'd29633: data = 8'h00;
      17'd29634: data = 8'hfe;
      17'd29635: data = 8'h00;
      17'd29636: data = 8'h00;
      17'd29637: data = 8'h02;
      17'd29638: data = 8'h04;
      17'd29639: data = 8'h04;
      17'd29640: data = 8'h04;
      17'd29641: data = 8'h04;
      17'd29642: data = 8'h05;
      17'd29643: data = 8'h06;
      17'd29644: data = 8'h04;
      17'd29645: data = 8'h04;
      17'd29646: data = 8'h02;
      17'd29647: data = 8'h01;
      17'd29648: data = 8'h00;
      17'd29649: data = 8'hfe;
      17'd29650: data = 8'h01;
      17'd29651: data = 8'h01;
      17'd29652: data = 8'h00;
      17'd29653: data = 8'h02;
      17'd29654: data = 8'h02;
      17'd29655: data = 8'h02;
      17'd29656: data = 8'h01;
      17'd29657: data = 8'h01;
      17'd29658: data = 8'h02;
      17'd29659: data = 8'h01;
      17'd29660: data = 8'h01;
      17'd29661: data = 8'h00;
      17'd29662: data = 8'hfe;
      17'd29663: data = 8'h00;
      17'd29664: data = 8'hfd;
      17'd29665: data = 8'hfe;
      17'd29666: data = 8'h00;
      17'd29667: data = 8'h00;
      17'd29668: data = 8'h01;
      17'd29669: data = 8'h02;
      17'd29670: data = 8'h04;
      17'd29671: data = 8'h02;
      17'd29672: data = 8'h01;
      17'd29673: data = 8'h02;
      17'd29674: data = 8'h02;
      17'd29675: data = 8'h00;
      17'd29676: data = 8'hfe;
      17'd29677: data = 8'hfe;
      17'd29678: data = 8'hfd;
      17'd29679: data = 8'hfd;
      17'd29680: data = 8'hfd;
      17'd29681: data = 8'hfe;
      17'd29682: data = 8'hfe;
      17'd29683: data = 8'hfe;
      17'd29684: data = 8'hfe;
      17'd29685: data = 8'h00;
      17'd29686: data = 8'h00;
      17'd29687: data = 8'h01;
      17'd29688: data = 8'h01;
      17'd29689: data = 8'h00;
      17'd29690: data = 8'hfd;
      17'd29691: data = 8'hfd;
      17'd29692: data = 8'hfd;
      17'd29693: data = 8'hfc;
      17'd29694: data = 8'hfc;
      17'd29695: data = 8'hfc;
      17'd29696: data = 8'hfc;
      17'd29697: data = 8'hfd;
      17'd29698: data = 8'hfd;
      17'd29699: data = 8'hfd;
      17'd29700: data = 8'hfe;
      17'd29701: data = 8'h01;
      17'd29702: data = 8'h00;
      17'd29703: data = 8'hfe;
      17'd29704: data = 8'h01;
      17'd29705: data = 8'h02;
      17'd29706: data = 8'h02;
      17'd29707: data = 8'h01;
      17'd29708: data = 8'h01;
      17'd29709: data = 8'h02;
      17'd29710: data = 8'h00;
      17'd29711: data = 8'h01;
      17'd29712: data = 8'h01;
      17'd29713: data = 8'h00;
      17'd29714: data = 8'h00;
      17'd29715: data = 8'h00;
      17'd29716: data = 8'h00;
      17'd29717: data = 8'hfe;
      17'd29718: data = 8'h00;
      17'd29719: data = 8'hfe;
      17'd29720: data = 8'hfe;
      17'd29721: data = 8'hfe;
      17'd29722: data = 8'h00;
      17'd29723: data = 8'h00;
      17'd29724: data = 8'h01;
      17'd29725: data = 8'h00;
      17'd29726: data = 8'hfe;
      17'd29727: data = 8'hfe;
      17'd29728: data = 8'hfe;
      17'd29729: data = 8'hfd;
      17'd29730: data = 8'hfa;
      17'd29731: data = 8'hfa;
      17'd29732: data = 8'hf9;
      17'd29733: data = 8'hf9;
      17'd29734: data = 8'hf9;
      17'd29735: data = 8'hfc;
      17'd29736: data = 8'hfd;
      17'd29737: data = 8'hfc;
      17'd29738: data = 8'hfd;
      17'd29739: data = 8'hfe;
      17'd29740: data = 8'hfd;
      17'd29741: data = 8'hfe;
      17'd29742: data = 8'hfe;
      17'd29743: data = 8'h00;
      17'd29744: data = 8'hfe;
      17'd29745: data = 8'hfd;
      17'd29746: data = 8'hfd;
      17'd29747: data = 8'hfd;
      17'd29748: data = 8'hfd;
      17'd29749: data = 8'hfd;
      17'd29750: data = 8'hfd;
      17'd29751: data = 8'hfd;
      17'd29752: data = 8'hfd;
      17'd29753: data = 8'hfe;
      17'd29754: data = 8'h00;
      17'd29755: data = 8'h00;
      17'd29756: data = 8'hfe;
      17'd29757: data = 8'hfd;
      17'd29758: data = 8'hfe;
      17'd29759: data = 8'hfd;
      17'd29760: data = 8'hfe;
      17'd29761: data = 8'hfd;
      17'd29762: data = 8'h00;
      17'd29763: data = 8'h00;
      17'd29764: data = 8'hfe;
      17'd29765: data = 8'hfc;
      17'd29766: data = 8'hfd;
      17'd29767: data = 8'hfd;
      17'd29768: data = 8'hfd;
      17'd29769: data = 8'hfe;
      17'd29770: data = 8'hfc;
      17'd29771: data = 8'hfd;
      17'd29772: data = 8'hfe;
      17'd29773: data = 8'hfe;
      17'd29774: data = 8'hfe;
      17'd29775: data = 8'h00;
      17'd29776: data = 8'h01;
      17'd29777: data = 8'h01;
      17'd29778: data = 8'hfe;
      17'd29779: data = 8'hfd;
      17'd29780: data = 8'hfe;
      17'd29781: data = 8'hfe;
      17'd29782: data = 8'hfe;
      17'd29783: data = 8'hfe;
      17'd29784: data = 8'hfe;
      17'd29785: data = 8'hfd;
      17'd29786: data = 8'hfe;
      17'd29787: data = 8'h00;
      17'd29788: data = 8'h00;
      17'd29789: data = 8'h00;
      17'd29790: data = 8'h00;
      17'd29791: data = 8'h00;
      17'd29792: data = 8'hfe;
      17'd29793: data = 8'hfd;
      17'd29794: data = 8'hfd;
      17'd29795: data = 8'hfe;
      17'd29796: data = 8'hfe;
      17'd29797: data = 8'hfe;
      17'd29798: data = 8'h01;
      17'd29799: data = 8'h01;
      17'd29800: data = 8'h00;
      17'd29801: data = 8'h01;
      17'd29802: data = 8'h01;
      17'd29803: data = 8'h01;
      17'd29804: data = 8'h01;
      17'd29805: data = 8'h00;
      17'd29806: data = 8'hfe;
      17'd29807: data = 8'h00;
      17'd29808: data = 8'hfe;
      17'd29809: data = 8'hfe;
      17'd29810: data = 8'hfd;
      17'd29811: data = 8'hfd;
      17'd29812: data = 8'hfd;
      17'd29813: data = 8'hfd;
      17'd29814: data = 8'hfe;
      17'd29815: data = 8'hfe;
      17'd29816: data = 8'hfe;
      17'd29817: data = 8'h00;
      17'd29818: data = 8'h01;
      17'd29819: data = 8'h00;
      17'd29820: data = 8'h00;
      17'd29821: data = 8'h00;
      17'd29822: data = 8'h00;
      17'd29823: data = 8'hfe;
      17'd29824: data = 8'hfd;
      17'd29825: data = 8'hfd;
      17'd29826: data = 8'hfd;
      17'd29827: data = 8'hfc;
      17'd29828: data = 8'hfd;
      17'd29829: data = 8'hfc;
      17'd29830: data = 8'hfd;
      17'd29831: data = 8'hfe;
      17'd29832: data = 8'h01;
      17'd29833: data = 8'h04;
      17'd29834: data = 8'h04;
      17'd29835: data = 8'h04;
      17'd29836: data = 8'h04;
      17'd29837: data = 8'h04;
      17'd29838: data = 8'h02;
      17'd29839: data = 8'h02;
      17'd29840: data = 8'hfe;
      17'd29841: data = 8'hfe;
      17'd29842: data = 8'hfd;
      17'd29843: data = 8'hfd;
      17'd29844: data = 8'hfd;
      17'd29845: data = 8'hfe;
      17'd29846: data = 8'h00;
      17'd29847: data = 8'h01;
      17'd29848: data = 8'h02;
      17'd29849: data = 8'h02;
      17'd29850: data = 8'h05;
      17'd29851: data = 8'h02;
      17'd29852: data = 8'h02;
      17'd29853: data = 8'h02;
      17'd29854: data = 8'h00;
      17'd29855: data = 8'hfd;
      17'd29856: data = 8'hfd;
      17'd29857: data = 8'hfa;
      17'd29858: data = 8'hf9;
      17'd29859: data = 8'hfc;
      17'd29860: data = 8'hfd;
      17'd29861: data = 8'h00;
      17'd29862: data = 8'h00;
      17'd29863: data = 8'h01;
      17'd29864: data = 8'h04;
      17'd29865: data = 8'h02;
      17'd29866: data = 8'h04;
      17'd29867: data = 8'h04;
      17'd29868: data = 8'h02;
      17'd29869: data = 8'h02;
      17'd29870: data = 8'h02;
      17'd29871: data = 8'h01;
      17'd29872: data = 8'h01;
      17'd29873: data = 8'h01;
      17'd29874: data = 8'h00;
      17'd29875: data = 8'h01;
      17'd29876: data = 8'h01;
      17'd29877: data = 8'h04;
      17'd29878: data = 8'h04;
      17'd29879: data = 8'h04;
      17'd29880: data = 8'h05;
      17'd29881: data = 8'h05;
      17'd29882: data = 8'h04;
      17'd29883: data = 8'h02;
      17'd29884: data = 8'h00;
      17'd29885: data = 8'hfd;
      17'd29886: data = 8'hfe;
      17'd29887: data = 8'h00;
      17'd29888: data = 8'h00;
      17'd29889: data = 8'h00;
      17'd29890: data = 8'h02;
      17'd29891: data = 8'h02;
      17'd29892: data = 8'h01;
      17'd29893: data = 8'h02;
      17'd29894: data = 8'h04;
      17'd29895: data = 8'h02;
      17'd29896: data = 8'h02;
      17'd29897: data = 8'h02;
      17'd29898: data = 8'h01;
      17'd29899: data = 8'h01;
      17'd29900: data = 8'h00;
      17'd29901: data = 8'hfe;
      17'd29902: data = 8'hfe;
      17'd29903: data = 8'h00;
      17'd29904: data = 8'h00;
      17'd29905: data = 8'h01;
      17'd29906: data = 8'h02;
      17'd29907: data = 8'h05;
      17'd29908: data = 8'h06;
      17'd29909: data = 8'h09;
      17'd29910: data = 8'h09;
      17'd29911: data = 8'h06;
      17'd29912: data = 8'h06;
      17'd29913: data = 8'h04;
      17'd29914: data = 8'h00;
      17'd29915: data = 8'hfd;
      17'd29916: data = 8'hfd;
      17'd29917: data = 8'hfe;
      17'd29918: data = 8'hfd;
      17'd29919: data = 8'h00;
      17'd29920: data = 8'hfe;
      17'd29921: data = 8'hfd;
      17'd29922: data = 8'hfe;
      17'd29923: data = 8'h01;
      17'd29924: data = 8'h02;
      17'd29925: data = 8'h02;
      17'd29926: data = 8'h01;
      17'd29927: data = 8'hfe;
      17'd29928: data = 8'hfd;
      17'd29929: data = 8'hfa;
      17'd29930: data = 8'hfa;
      17'd29931: data = 8'hf9;
      17'd29932: data = 8'hf9;
      17'd29933: data = 8'hfc;
      17'd29934: data = 8'hfa;
      17'd29935: data = 8'hfc;
      17'd29936: data = 8'hfe;
      17'd29937: data = 8'hfe;
      17'd29938: data = 8'h00;
      17'd29939: data = 8'h01;
      17'd29940: data = 8'h00;
      17'd29941: data = 8'h01;
      17'd29942: data = 8'h02;
      17'd29943: data = 8'h01;
      17'd29944: data = 8'h00;
      17'd29945: data = 8'hfe;
      17'd29946: data = 8'h00;
      17'd29947: data = 8'h01;
      17'd29948: data = 8'h01;
      17'd29949: data = 8'h00;
      17'd29950: data = 8'h01;
      17'd29951: data = 8'h01;
      17'd29952: data = 8'h02;
      17'd29953: data = 8'h02;
      17'd29954: data = 8'h02;
      17'd29955: data = 8'h02;
      17'd29956: data = 8'h01;
      17'd29957: data = 8'h01;
      17'd29958: data = 8'h00;
      17'd29959: data = 8'hfe;
      17'd29960: data = 8'hfd;
      17'd29961: data = 8'hfd;
      17'd29962: data = 8'hfe;
      17'd29963: data = 8'hfc;
      17'd29964: data = 8'hfc;
      17'd29965: data = 8'hfd;
      17'd29966: data = 8'hfd;
      17'd29967: data = 8'hfd;
      17'd29968: data = 8'hfc;
      17'd29969: data = 8'hfc;
      17'd29970: data = 8'hfd;
      17'd29971: data = 8'hfc;
      17'd29972: data = 8'hf9;
      17'd29973: data = 8'hfa;
      17'd29974: data = 8'hfa;
      17'd29975: data = 8'hfa;
      17'd29976: data = 8'hf9;
      17'd29977: data = 8'hfa;
      17'd29978: data = 8'hf9;
      17'd29979: data = 8'hfc;
      17'd29980: data = 8'hfa;
      17'd29981: data = 8'hfc;
      17'd29982: data = 8'hfd;
      17'd29983: data = 8'hfe;
      17'd29984: data = 8'hfe;
      17'd29985: data = 8'hfe;
      17'd29986: data = 8'hfe;
      17'd29987: data = 8'hfc;
      17'd29988: data = 8'hfc;
      17'd29989: data = 8'hfa;
      17'd29990: data = 8'hfa;
      17'd29991: data = 8'hfc;
      17'd29992: data = 8'hfc;
      17'd29993: data = 8'hfa;
      17'd29994: data = 8'hfd;
      17'd29995: data = 8'hfe;
      17'd29996: data = 8'h00;
      17'd29997: data = 8'h00;
      17'd29998: data = 8'h00;
      17'd29999: data = 8'h00;
      17'd30000: data = 8'hfe;
      17'd30001: data = 8'h01;
      17'd30002: data = 8'hfe;
      17'd30003: data = 8'hfc;
      17'd30004: data = 8'hfd;
      17'd30005: data = 8'hfc;
      17'd30006: data = 8'hfd;
      17'd30007: data = 8'hfe;
      17'd30008: data = 8'hfe;
      17'd30009: data = 8'hfe;
      17'd30010: data = 8'h01;
      17'd30011: data = 8'h00;
      17'd30012: data = 8'h01;
      17'd30013: data = 8'h01;
      17'd30014: data = 8'h00;
      17'd30015: data = 8'h01;
      17'd30016: data = 8'hfd;
      17'd30017: data = 8'hfd;
      17'd30018: data = 8'hfc;
      17'd30019: data = 8'hfa;
      17'd30020: data = 8'hf9;
      17'd30021: data = 8'hfa;
      17'd30022: data = 8'hf9;
      17'd30023: data = 8'hfc;
      17'd30024: data = 8'hfe;
      17'd30025: data = 8'hfd;
      17'd30026: data = 8'h00;
      17'd30027: data = 8'h01;
      17'd30028: data = 8'h00;
      17'd30029: data = 8'hfe;
      17'd30030: data = 8'hfd;
      17'd30031: data = 8'hfd;
      17'd30032: data = 8'hfd;
      17'd30033: data = 8'hfd;
      17'd30034: data = 8'hfc;
      17'd30035: data = 8'hfc;
      17'd30036: data = 8'hfe;
      17'd30037: data = 8'h00;
      17'd30038: data = 8'h01;
      17'd30039: data = 8'h01;
      17'd30040: data = 8'h01;
      17'd30041: data = 8'h01;
      17'd30042: data = 8'h02;
      17'd30043: data = 8'h02;
      17'd30044: data = 8'h01;
      17'd30045: data = 8'h00;
      17'd30046: data = 8'hfd;
      17'd30047: data = 8'hfd;
      17'd30048: data = 8'hfc;
      17'd30049: data = 8'hfc;
      17'd30050: data = 8'hfc;
      17'd30051: data = 8'hfe;
      17'd30052: data = 8'h00;
      17'd30053: data = 8'hfe;
      17'd30054: data = 8'h00;
      17'd30055: data = 8'h01;
      17'd30056: data = 8'h00;
      17'd30057: data = 8'h02;
      17'd30058: data = 8'h02;
      17'd30059: data = 8'h00;
      17'd30060: data = 8'hfe;
      17'd30061: data = 8'hfd;
      17'd30062: data = 8'hfc;
      17'd30063: data = 8'hfc;
      17'd30064: data = 8'hfa;
      17'd30065: data = 8'hf9;
      17'd30066: data = 8'hfc;
      17'd30067: data = 8'hfd;
      17'd30068: data = 8'hfe;
      17'd30069: data = 8'h02;
      17'd30070: data = 8'h02;
      17'd30071: data = 8'h04;
      17'd30072: data = 8'h05;
      17'd30073: data = 8'h04;
      17'd30074: data = 8'h01;
      17'd30075: data = 8'h00;
      17'd30076: data = 8'hfe;
      17'd30077: data = 8'hfe;
      17'd30078: data = 8'h00;
      17'd30079: data = 8'hfe;
      17'd30080: data = 8'hfd;
      17'd30081: data = 8'h00;
      17'd30082: data = 8'h01;
      17'd30083: data = 8'h01;
      17'd30084: data = 8'h02;
      17'd30085: data = 8'h05;
      17'd30086: data = 8'h04;
      17'd30087: data = 8'h04;
      17'd30088: data = 8'h04;
      17'd30089: data = 8'h02;
      17'd30090: data = 8'h01;
      17'd30091: data = 8'h00;
      17'd30092: data = 8'hfd;
      17'd30093: data = 8'hfc;
      17'd30094: data = 8'hfc;
      17'd30095: data = 8'hfd;
      17'd30096: data = 8'hfd;
      17'd30097: data = 8'hfd;
      17'd30098: data = 8'h00;
      17'd30099: data = 8'h00;
      17'd30100: data = 8'h00;
      17'd30101: data = 8'h02;
      17'd30102: data = 8'h02;
      17'd30103: data = 8'h01;
      17'd30104: data = 8'h01;
      17'd30105: data = 8'h00;
      17'd30106: data = 8'hfe;
      17'd30107: data = 8'h00;
      17'd30108: data = 8'hfe;
      17'd30109: data = 8'hfd;
      17'd30110: data = 8'hfe;
      17'd30111: data = 8'hfe;
      17'd30112: data = 8'h00;
      17'd30113: data = 8'h01;
      17'd30114: data = 8'h02;
      17'd30115: data = 8'h05;
      17'd30116: data = 8'h05;
      17'd30117: data = 8'h05;
      17'd30118: data = 8'h06;
      17'd30119: data = 8'h04;
      17'd30120: data = 8'h02;
      17'd30121: data = 8'h02;
      17'd30122: data = 8'h00;
      17'd30123: data = 8'h00;
      17'd30124: data = 8'hfe;
      17'd30125: data = 8'h00;
      17'd30126: data = 8'h01;
      17'd30127: data = 8'h00;
      17'd30128: data = 8'h01;
      17'd30129: data = 8'h04;
      17'd30130: data = 8'h04;
      17'd30131: data = 8'h04;
      17'd30132: data = 8'h04;
      17'd30133: data = 8'h02;
      17'd30134: data = 8'h02;
      17'd30135: data = 8'h01;
      17'd30136: data = 8'h01;
      17'd30137: data = 8'hfe;
      17'd30138: data = 8'hfd;
      17'd30139: data = 8'h00;
      17'd30140: data = 8'h00;
      17'd30141: data = 8'hfe;
      17'd30142: data = 8'h02;
      17'd30143: data = 8'h04;
      17'd30144: data = 8'h04;
      17'd30145: data = 8'h05;
      17'd30146: data = 8'h05;
      17'd30147: data = 8'h05;
      17'd30148: data = 8'h04;
      17'd30149: data = 8'h02;
      17'd30150: data = 8'h01;
      17'd30151: data = 8'h00;
      17'd30152: data = 8'hfe;
      17'd30153: data = 8'hfa;
      17'd30154: data = 8'hfc;
      17'd30155: data = 8'hfc;
      17'd30156: data = 8'hf9;
      17'd30157: data = 8'hfa;
      17'd30158: data = 8'hfc;
      17'd30159: data = 8'hfd;
      17'd30160: data = 8'hfe;
      17'd30161: data = 8'h00;
      17'd30162: data = 8'h00;
      17'd30163: data = 8'hfe;
      17'd30164: data = 8'hfd;
      17'd30165: data = 8'hfc;
      17'd30166: data = 8'hfc;
      17'd30167: data = 8'hfa;
      17'd30168: data = 8'hf9;
      17'd30169: data = 8'hf9;
      17'd30170: data = 8'hfa;
      17'd30171: data = 8'hfa;
      17'd30172: data = 8'hfc;
      17'd30173: data = 8'hfe;
      17'd30174: data = 8'h00;
      17'd30175: data = 8'h00;
      17'd30176: data = 8'h01;
      17'd30177: data = 8'h04;
      17'd30178: data = 8'h02;
      17'd30179: data = 8'h02;
      17'd30180: data = 8'h04;
      17'd30181: data = 8'h02;
      17'd30182: data = 8'h01;
      17'd30183: data = 8'h01;
      17'd30184: data = 8'h01;
      17'd30185: data = 8'h02;
      17'd30186: data = 8'h01;
      17'd30187: data = 8'h01;
      17'd30188: data = 8'h01;
      17'd30189: data = 8'h04;
      17'd30190: data = 8'h05;
      17'd30191: data = 8'h05;
      17'd30192: data = 8'h04;
      17'd30193: data = 8'h02;
      17'd30194: data = 8'h02;
      17'd30195: data = 8'h01;
      17'd30196: data = 8'h00;
      17'd30197: data = 8'hfe;
      17'd30198: data = 8'hfc;
      17'd30199: data = 8'hfc;
      17'd30200: data = 8'hfc;
      17'd30201: data = 8'hfa;
      17'd30202: data = 8'hf9;
      17'd30203: data = 8'hfa;
      17'd30204: data = 8'hfa;
      17'd30205: data = 8'hfa;
      17'd30206: data = 8'hfa;
      17'd30207: data = 8'hfa;
      17'd30208: data = 8'hfa;
      17'd30209: data = 8'hfc;
      17'd30210: data = 8'hfc;
      17'd30211: data = 8'hfc;
      17'd30212: data = 8'hfa;
      17'd30213: data = 8'hf9;
      17'd30214: data = 8'hfa;
      17'd30215: data = 8'hf9;
      17'd30216: data = 8'hfa;
      17'd30217: data = 8'hfa;
      17'd30218: data = 8'hfc;
      17'd30219: data = 8'hfd;
      17'd30220: data = 8'h00;
      17'd30221: data = 8'h00;
      17'd30222: data = 8'hfe;
      17'd30223: data = 8'h01;
      17'd30224: data = 8'h01;
      17'd30225: data = 8'h01;
      17'd30226: data = 8'hfe;
      17'd30227: data = 8'hfe;
      17'd30228: data = 8'hfe;
      17'd30229: data = 8'h00;
      17'd30230: data = 8'hfe;
      17'd30231: data = 8'h01;
      17'd30232: data = 8'h02;
      17'd30233: data = 8'h04;
      17'd30234: data = 8'h04;
      17'd30235: data = 8'h04;
      17'd30236: data = 8'h04;
      17'd30237: data = 8'h04;
      17'd30238: data = 8'h04;
      17'd30239: data = 8'h02;
      17'd30240: data = 8'h00;
      17'd30241: data = 8'h00;
      17'd30242: data = 8'h00;
      17'd30243: data = 8'hfd;
      17'd30244: data = 8'hfd;
      17'd30245: data = 8'hfd;
      17'd30246: data = 8'hfe;
      17'd30247: data = 8'hfd;
      17'd30248: data = 8'hfd;
      17'd30249: data = 8'hfe;
      17'd30250: data = 8'hfe;
      17'd30251: data = 8'hfe;
      17'd30252: data = 8'hfe;
      17'd30253: data = 8'hfc;
      17'd30254: data = 8'hfc;
      17'd30255: data = 8'hfa;
      17'd30256: data = 8'hfa;
      17'd30257: data = 8'hf9;
      17'd30258: data = 8'hf6;
      17'd30259: data = 8'hf6;
      17'd30260: data = 8'hf9;
      17'd30261: data = 8'hf9;
      17'd30262: data = 8'hf9;
      17'd30263: data = 8'hfa;
      17'd30264: data = 8'hfa;
      17'd30265: data = 8'hfc;
      17'd30266: data = 8'hfd;
      17'd30267: data = 8'hfd;
      17'd30268: data = 8'hfe;
      17'd30269: data = 8'hfd;
      17'd30270: data = 8'hfe;
      17'd30271: data = 8'hfe;
      17'd30272: data = 8'h00;
      17'd30273: data = 8'hfe;
      17'd30274: data = 8'hfe;
      17'd30275: data = 8'h00;
      17'd30276: data = 8'h01;
      17'd30277: data = 8'h01;
      17'd30278: data = 8'h00;
      17'd30279: data = 8'h01;
      17'd30280: data = 8'h02;
      17'd30281: data = 8'h02;
      17'd30282: data = 8'h02;
      17'd30283: data = 8'h01;
      17'd30284: data = 8'h01;
      17'd30285: data = 8'h01;
      17'd30286: data = 8'h01;
      17'd30287: data = 8'h00;
      17'd30288: data = 8'h00;
      17'd30289: data = 8'h00;
      17'd30290: data = 8'h00;
      17'd30291: data = 8'h01;
      17'd30292: data = 8'h01;
      17'd30293: data = 8'h01;
      17'd30294: data = 8'h01;
      17'd30295: data = 8'h01;
      17'd30296: data = 8'h01;
      17'd30297: data = 8'hfe;
      17'd30298: data = 8'hfd;
      17'd30299: data = 8'hfd;
      17'd30300: data = 8'hf9;
      17'd30301: data = 8'hfa;
      17'd30302: data = 8'hfa;
      17'd30303: data = 8'hf9;
      17'd30304: data = 8'hfa;
      17'd30305: data = 8'hfa;
      17'd30306: data = 8'hf9;
      17'd30307: data = 8'hfc;
      17'd30308: data = 8'hfd;
      17'd30309: data = 8'hfd;
      17'd30310: data = 8'hfd;
      17'd30311: data = 8'hfd;
      17'd30312: data = 8'hfd;
      17'd30313: data = 8'hfc;
      17'd30314: data = 8'hfc;
      17'd30315: data = 8'hfc;
      17'd30316: data = 8'hfc;
      17'd30317: data = 8'hfc;
      17'd30318: data = 8'hfd;
      17'd30319: data = 8'hfe;
      17'd30320: data = 8'h01;
      17'd30321: data = 8'h01;
      17'd30322: data = 8'h00;
      17'd30323: data = 8'h02;
      17'd30324: data = 8'h02;
      17'd30325: data = 8'h02;
      17'd30326: data = 8'h04;
      17'd30327: data = 8'h02;
      17'd30328: data = 8'h00;
      17'd30329: data = 8'h01;
      17'd30330: data = 8'h01;
      17'd30331: data = 8'h01;
      17'd30332: data = 8'h02;
      17'd30333: data = 8'h01;
      17'd30334: data = 8'h02;
      17'd30335: data = 8'h04;
      17'd30336: data = 8'h01;
      17'd30337: data = 8'h01;
      17'd30338: data = 8'h04;
      17'd30339: data = 8'h01;
      17'd30340: data = 8'h01;
      17'd30341: data = 8'h02;
      17'd30342: data = 8'h01;
      17'd30343: data = 8'h00;
      17'd30344: data = 8'h01;
      17'd30345: data = 8'h02;
      17'd30346: data = 8'h01;
      17'd30347: data = 8'h00;
      17'd30348: data = 8'h01;
      17'd30349: data = 8'h01;
      17'd30350: data = 8'h00;
      17'd30351: data = 8'h00;
      17'd30352: data = 8'h00;
      17'd30353: data = 8'h01;
      17'd30354: data = 8'h00;
      17'd30355: data = 8'h00;
      17'd30356: data = 8'h00;
      17'd30357: data = 8'hfe;
      17'd30358: data = 8'hfe;
      17'd30359: data = 8'h00;
      17'd30360: data = 8'hfe;
      17'd30361: data = 8'hfc;
      17'd30362: data = 8'hfe;
      17'd30363: data = 8'hfe;
      17'd30364: data = 8'hfe;
      17'd30365: data = 8'h00;
      17'd30366: data = 8'h00;
      17'd30367: data = 8'h00;
      17'd30368: data = 8'h01;
      17'd30369: data = 8'h00;
      17'd30370: data = 8'h01;
      17'd30371: data = 8'h02;
      17'd30372: data = 8'h02;
      17'd30373: data = 8'h01;
      17'd30374: data = 8'h01;
      17'd30375: data = 8'h02;
      17'd30376: data = 8'h02;
      17'd30377: data = 8'h02;
      17'd30378: data = 8'h04;
      17'd30379: data = 8'h05;
      17'd30380: data = 8'h05;
      17'd30381: data = 8'h06;
      17'd30382: data = 8'h09;
      17'd30383: data = 8'h09;
      17'd30384: data = 8'h0a;
      17'd30385: data = 8'h0a;
      17'd30386: data = 8'h06;
      17'd30387: data = 8'h05;
      17'd30388: data = 8'h04;
      17'd30389: data = 8'h02;
      17'd30390: data = 8'h01;
      17'd30391: data = 8'h01;
      17'd30392: data = 8'h01;
      17'd30393: data = 8'h01;
      17'd30394: data = 8'h00;
      17'd30395: data = 8'h00;
      17'd30396: data = 8'h00;
      17'd30397: data = 8'hfe;
      17'd30398: data = 8'hfd;
      17'd30399: data = 8'hfd;
      17'd30400: data = 8'hfc;
      17'd30401: data = 8'hfa;
      17'd30402: data = 8'hfa;
      17'd30403: data = 8'hf9;
      17'd30404: data = 8'hfa;
      17'd30405: data = 8'hfa;
      17'd30406: data = 8'hf9;
      17'd30407: data = 8'hfa;
      17'd30408: data = 8'hf9;
      17'd30409: data = 8'hf9;
      17'd30410: data = 8'hf6;
      17'd30411: data = 8'hf6;
      17'd30412: data = 8'hfc;
      17'd30413: data = 8'hfc;
      17'd30414: data = 8'hfc;
      17'd30415: data = 8'hfd;
      17'd30416: data = 8'hfe;
      17'd30417: data = 8'h00;
      17'd30418: data = 8'h00;
      17'd30419: data = 8'h00;
      17'd30420: data = 8'h00;
      17'd30421: data = 8'h02;
      17'd30422: data = 8'h04;
      17'd30423: data = 8'h04;
      17'd30424: data = 8'h05;
      17'd30425: data = 8'h04;
      17'd30426: data = 8'h05;
      17'd30427: data = 8'h04;
      17'd30428: data = 8'h02;
      17'd30429: data = 8'h05;
      17'd30430: data = 8'h05;
      17'd30431: data = 8'h06;
      17'd30432: data = 8'h09;
      17'd30433: data = 8'h06;
      17'd30434: data = 8'h05;
      17'd30435: data = 8'h05;
      17'd30436: data = 8'h05;
      17'd30437: data = 8'h04;
      17'd30438: data = 8'h02;
      17'd30439: data = 8'h02;
      17'd30440: data = 8'h02;
      17'd30441: data = 8'h00;
      17'd30442: data = 8'hfe;
      17'd30443: data = 8'hfe;
      17'd30444: data = 8'hfd;
      17'd30445: data = 8'hfc;
      17'd30446: data = 8'hfd;
      17'd30447: data = 8'hfc;
      17'd30448: data = 8'hfa;
      17'd30449: data = 8'hfc;
      17'd30450: data = 8'hfa;
      17'd30451: data = 8'hf9;
      17'd30452: data = 8'hfa;
      17'd30453: data = 8'hfa;
      17'd30454: data = 8'hfa;
      17'd30455: data = 8'hfa;
      17'd30456: data = 8'hfa;
      17'd30457: data = 8'hfa;
      17'd30458: data = 8'hf9;
      17'd30459: data = 8'hf6;
      17'd30460: data = 8'hf9;
      17'd30461: data = 8'hf6;
      17'd30462: data = 8'hfa;
      17'd30463: data = 8'hfa;
      17'd30464: data = 8'hfa;
      17'd30465: data = 8'hfd;
      17'd30466: data = 8'hfd;
      17'd30467: data = 8'hfe;
      17'd30468: data = 8'h00;
      17'd30469: data = 8'h01;
      17'd30470: data = 8'h01;
      17'd30471: data = 8'hfe;
      17'd30472: data = 8'h02;
      17'd30473: data = 8'h04;
      17'd30474: data = 8'h02;
      17'd30475: data = 8'h02;
      17'd30476: data = 8'h02;
      17'd30477: data = 8'h04;
      17'd30478: data = 8'h04;
      17'd30479: data = 8'h04;
      17'd30480: data = 8'h05;
      17'd30481: data = 8'h04;
      17'd30482: data = 8'h05;
      17'd30483: data = 8'h05;
      17'd30484: data = 8'h06;
      17'd30485: data = 8'h05;
      17'd30486: data = 8'h04;
      17'd30487: data = 8'h04;
      17'd30488: data = 8'h01;
      17'd30489: data = 8'h00;
      17'd30490: data = 8'h00;
      17'd30491: data = 8'h00;
      17'd30492: data = 8'hfd;
      17'd30493: data = 8'hfd;
      17'd30494: data = 8'hfd;
      17'd30495: data = 8'hfd;
      17'd30496: data = 8'hfd;
      17'd30497: data = 8'hfd;
      17'd30498: data = 8'hfe;
      17'd30499: data = 8'hfe;
      17'd30500: data = 8'hfd;
      17'd30501: data = 8'hf9;
      17'd30502: data = 8'hf9;
      17'd30503: data = 8'hf9;
      17'd30504: data = 8'hf6;
      17'd30505: data = 8'hf5;
      17'd30506: data = 8'hf6;
      17'd30507: data = 8'hf6;
      17'd30508: data = 8'hfa;
      17'd30509: data = 8'hfc;
      17'd30510: data = 8'hfd;
      17'd30511: data = 8'hfd;
      17'd30512: data = 8'hfe;
      17'd30513: data = 8'h00;
      17'd30514: data = 8'hfe;
      17'd30515: data = 8'hfd;
      17'd30516: data = 8'hfd;
      17'd30517: data = 8'hfd;
      17'd30518: data = 8'hfd;
      17'd30519: data = 8'hfd;
      17'd30520: data = 8'hfc;
      17'd30521: data = 8'hfd;
      17'd30522: data = 8'hfe;
      17'd30523: data = 8'h00;
      17'd30524: data = 8'h02;
      17'd30525: data = 8'h01;
      17'd30526: data = 8'h04;
      17'd30527: data = 8'h05;
      17'd30528: data = 8'h06;
      17'd30529: data = 8'h06;
      17'd30530: data = 8'h05;
      17'd30531: data = 8'h06;
      17'd30532: data = 8'h02;
      17'd30533: data = 8'h04;
      17'd30534: data = 8'h02;
      17'd30535: data = 8'h00;
      17'd30536: data = 8'h00;
      17'd30537: data = 8'hfe;
      17'd30538: data = 8'hfe;
      17'd30539: data = 8'hfe;
      17'd30540: data = 8'h01;
      17'd30541: data = 8'h02;
      17'd30542: data = 8'h04;
      17'd30543: data = 8'h04;
      17'd30544: data = 8'h04;
      17'd30545: data = 8'h02;
      17'd30546: data = 8'h01;
      17'd30547: data = 8'h00;
      17'd30548: data = 8'hfe;
      17'd30549: data = 8'hfd;
      17'd30550: data = 8'hfd;
      17'd30551: data = 8'hfc;
      17'd30552: data = 8'hfa;
      17'd30553: data = 8'hfa;
      17'd30554: data = 8'hfa;
      17'd30555: data = 8'hfc;
      17'd30556: data = 8'hfe;
      17'd30557: data = 8'hfd;
      17'd30558: data = 8'hfe;
      17'd30559: data = 8'hfe;
      17'd30560: data = 8'h00;
      17'd30561: data = 8'hfe;
      17'd30562: data = 8'hfd;
      17'd30563: data = 8'hfc;
      17'd30564: data = 8'hfa;
      17'd30565: data = 8'hfa;
      17'd30566: data = 8'hfa;
      17'd30567: data = 8'hfc;
      17'd30568: data = 8'hfc;
      17'd30569: data = 8'hfd;
      17'd30570: data = 8'hfe;
      17'd30571: data = 8'h00;
      17'd30572: data = 8'h01;
      17'd30573: data = 8'h01;
      17'd30574: data = 8'h02;
      17'd30575: data = 8'h02;
      17'd30576: data = 8'h04;
      17'd30577: data = 8'h02;
      17'd30578: data = 8'h04;
      17'd30579: data = 8'h02;
      17'd30580: data = 8'h01;
      17'd30581: data = 8'h01;
      17'd30582: data = 8'h01;
      17'd30583: data = 8'h01;
      17'd30584: data = 8'h02;
      17'd30585: data = 8'h02;
      17'd30586: data = 8'h04;
      17'd30587: data = 8'h05;
      17'd30588: data = 8'h05;
      17'd30589: data = 8'h04;
      17'd30590: data = 8'h05;
      17'd30591: data = 8'h05;
      17'd30592: data = 8'h02;
      17'd30593: data = 8'h01;
      17'd30594: data = 8'hfe;
      17'd30595: data = 8'hfd;
      17'd30596: data = 8'hfc;
      17'd30597: data = 8'hfa;
      17'd30598: data = 8'hfa;
      17'd30599: data = 8'hfa;
      17'd30600: data = 8'hfa;
      17'd30601: data = 8'hfd;
      17'd30602: data = 8'hfd;
      17'd30603: data = 8'h00;
      17'd30604: data = 8'h01;
      17'd30605: data = 8'h00;
      17'd30606: data = 8'hfd;
      17'd30607: data = 8'hfd;
      17'd30608: data = 8'hfd;
      17'd30609: data = 8'hfc;
      17'd30610: data = 8'hfc;
      17'd30611: data = 8'hfc;
      17'd30612: data = 8'hfd;
      17'd30613: data = 8'hfc;
      17'd30614: data = 8'hfe;
      17'd30615: data = 8'h01;
      17'd30616: data = 8'h02;
      17'd30617: data = 8'h05;
      17'd30618: data = 8'h06;
      17'd30619: data = 8'h09;
      17'd30620: data = 8'h06;
      17'd30621: data = 8'h05;
      17'd30622: data = 8'h05;
      17'd30623: data = 8'h05;
      17'd30624: data = 8'h01;
      17'd30625: data = 8'h02;
      17'd30626: data = 8'h00;
      17'd30627: data = 8'h01;
      17'd30628: data = 8'h01;
      17'd30629: data = 8'h01;
      17'd30630: data = 8'h02;
      17'd30631: data = 8'h02;
      17'd30632: data = 8'h04;
      17'd30633: data = 8'h04;
      17'd30634: data = 8'h02;
      17'd30635: data = 8'h01;
      17'd30636: data = 8'h00;
      17'd30637: data = 8'h00;
      17'd30638: data = 8'h00;
      17'd30639: data = 8'hfd;
      17'd30640: data = 8'hfd;
      17'd30641: data = 8'hfa;
      17'd30642: data = 8'hfa;
      17'd30643: data = 8'hfa;
      17'd30644: data = 8'hfa;
      17'd30645: data = 8'hf9;
      17'd30646: data = 8'hfa;
      17'd30647: data = 8'hfc;
      17'd30648: data = 8'hfd;
      17'd30649: data = 8'hfd;
      17'd30650: data = 8'hfd;
      17'd30651: data = 8'hfe;
      17'd30652: data = 8'hfe;
      17'd30653: data = 8'hfe;
      17'd30654: data = 8'hfe;
      17'd30655: data = 8'hfe;
      17'd30656: data = 8'hfd;
      17'd30657: data = 8'hfd;
      17'd30658: data = 8'hfe;
      17'd30659: data = 8'hfe;
      17'd30660: data = 8'hfe;
      17'd30661: data = 8'h01;
      17'd30662: data = 8'h01;
      17'd30663: data = 8'h01;
      17'd30664: data = 8'h01;
      17'd30665: data = 8'h02;
      17'd30666: data = 8'h02;
      17'd30667: data = 8'h02;
      17'd30668: data = 8'h02;
      17'd30669: data = 8'h02;
      17'd30670: data = 8'h02;
      17'd30671: data = 8'h02;
      17'd30672: data = 8'h02;
      17'd30673: data = 8'h02;
      17'd30674: data = 8'h02;
      17'd30675: data = 8'h01;
      17'd30676: data = 8'hfe;
      17'd30677: data = 8'h00;
      17'd30678: data = 8'h00;
      17'd30679: data = 8'hfe;
      17'd30680: data = 8'h00;
      17'd30681: data = 8'h00;
      17'd30682: data = 8'hfd;
      17'd30683: data = 8'hfe;
      17'd30684: data = 8'hfe;
      17'd30685: data = 8'hfd;
      17'd30686: data = 8'hfd;
      17'd30687: data = 8'hfd;
      17'd30688: data = 8'hfd;
      17'd30689: data = 8'hfd;
      17'd30690: data = 8'hfd;
      17'd30691: data = 8'hfc;
      17'd30692: data = 8'hfc;
      17'd30693: data = 8'hfc;
      17'd30694: data = 8'hfc;
      17'd30695: data = 8'hfc;
      17'd30696: data = 8'hfa;
      17'd30697: data = 8'hfa;
      17'd30698: data = 8'hf9;
      17'd30699: data = 8'hfa;
      17'd30700: data = 8'hf9;
      17'd30701: data = 8'hfa;
      17'd30702: data = 8'hfa;
      17'd30703: data = 8'hfc;
      17'd30704: data = 8'hfa;
      17'd30705: data = 8'hfa;
      17'd30706: data = 8'hfd;
      17'd30707: data = 8'hfd;
      17'd30708: data = 8'h00;
      17'd30709: data = 8'h00;
      17'd30710: data = 8'h00;
      17'd30711: data = 8'h01;
      17'd30712: data = 8'h00;
      17'd30713: data = 8'hfe;
      17'd30714: data = 8'h01;
      17'd30715: data = 8'h01;
      17'd30716: data = 8'h01;
      17'd30717: data = 8'h02;
      17'd30718: data = 8'h02;
      17'd30719: data = 8'h01;
      17'd30720: data = 8'h02;
      17'd30721: data = 8'h02;
      17'd30722: data = 8'h02;
      17'd30723: data = 8'h02;
      17'd30724: data = 8'h01;
      17'd30725: data = 8'h01;
      17'd30726: data = 8'h00;
      17'd30727: data = 8'h00;
      17'd30728: data = 8'h00;
      17'd30729: data = 8'h00;
      17'd30730: data = 8'h00;
      17'd30731: data = 8'hfe;
      17'd30732: data = 8'hfd;
      17'd30733: data = 8'hfe;
      17'd30734: data = 8'hfe;
      17'd30735: data = 8'hfe;
      17'd30736: data = 8'h00;
      17'd30737: data = 8'hfe;
      17'd30738: data = 8'hfe;
      17'd30739: data = 8'hfd;
      17'd30740: data = 8'hfa;
      17'd30741: data = 8'hfa;
      17'd30742: data = 8'hfc;
      17'd30743: data = 8'hfa;
      17'd30744: data = 8'hf9;
      17'd30745: data = 8'hfc;
      17'd30746: data = 8'hfc;
      17'd30747: data = 8'hfd;
      17'd30748: data = 8'hfe;
      17'd30749: data = 8'hfd;
      17'd30750: data = 8'hfe;
      17'd30751: data = 8'hfd;
      17'd30752: data = 8'hfc;
      17'd30753: data = 8'hfe;
      17'd30754: data = 8'hfe;
      17'd30755: data = 8'hfe;
      17'd30756: data = 8'hfe;
      17'd30757: data = 8'hfe;
      17'd30758: data = 8'hfe;
      17'd30759: data = 8'hfe;
      17'd30760: data = 8'hfd;
      17'd30761: data = 8'h00;
      17'd30762: data = 8'h00;
      17'd30763: data = 8'h01;
      17'd30764: data = 8'h02;
      17'd30765: data = 8'h02;
      17'd30766: data = 8'h04;
      17'd30767: data = 8'h01;
      17'd30768: data = 8'h01;
      17'd30769: data = 8'h01;
      17'd30770: data = 8'h01;
      17'd30771: data = 8'h01;
      17'd30772: data = 8'h01;
      17'd30773: data = 8'h00;
      17'd30774: data = 8'h00;
      17'd30775: data = 8'h01;
      17'd30776: data = 8'h01;
      17'd30777: data = 8'h00;
      17'd30778: data = 8'h01;
      17'd30779: data = 8'h02;
      17'd30780: data = 8'h04;
      17'd30781: data = 8'h02;
      17'd30782: data = 8'h02;
      17'd30783: data = 8'h01;
      17'd30784: data = 8'h00;
      17'd30785: data = 8'h00;
      17'd30786: data = 8'hfe;
      17'd30787: data = 8'hfe;
      17'd30788: data = 8'hfe;
      17'd30789: data = 8'hfd;
      17'd30790: data = 8'hfe;
      17'd30791: data = 8'hfd;
      17'd30792: data = 8'hfd;
      17'd30793: data = 8'hfe;
      17'd30794: data = 8'h00;
      17'd30795: data = 8'hfe;
      17'd30796: data = 8'hfd;
      17'd30797: data = 8'hfd;
      17'd30798: data = 8'hfc;
      17'd30799: data = 8'hfc;
      17'd30800: data = 8'hfc;
      17'd30801: data = 8'hfc;
      17'd30802: data = 8'hfd;
      17'd30803: data = 8'hfe;
      17'd30804: data = 8'hfd;
      17'd30805: data = 8'hfd;
      17'd30806: data = 8'hfd;
      17'd30807: data = 8'hfe;
      17'd30808: data = 8'hfd;
      17'd30809: data = 8'h00;
      17'd30810: data = 8'h00;
      17'd30811: data = 8'h01;
      17'd30812: data = 8'hfe;
      17'd30813: data = 8'hfd;
      17'd30814: data = 8'h02;
      17'd30815: data = 8'hfe;
      17'd30816: data = 8'h00;
      17'd30817: data = 8'h01;
      17'd30818: data = 8'h01;
      17'd30819: data = 8'h02;
      17'd30820: data = 8'h04;
      17'd30821: data = 8'h02;
      17'd30822: data = 8'h04;
      17'd30823: data = 8'h02;
      17'd30824: data = 8'h02;
      17'd30825: data = 8'h02;
      17'd30826: data = 8'h01;
      17'd30827: data = 8'h02;
      17'd30828: data = 8'h01;
      17'd30829: data = 8'h00;
      17'd30830: data = 8'h00;
      17'd30831: data = 8'h00;
      17'd30832: data = 8'hfe;
      17'd30833: data = 8'hfd;
      17'd30834: data = 8'hfe;
      17'd30835: data = 8'hfe;
      17'd30836: data = 8'hfe;
      17'd30837: data = 8'hfe;
      17'd30838: data = 8'hfe;
      17'd30839: data = 8'h00;
      17'd30840: data = 8'h00;
      17'd30841: data = 8'hfe;
      17'd30842: data = 8'hfe;
      17'd30843: data = 8'hfe;
      17'd30844: data = 8'hfe;
      17'd30845: data = 8'hfe;
      17'd30846: data = 8'hfe;
      17'd30847: data = 8'h01;
      17'd30848: data = 8'hf6;
      17'd30849: data = 8'hfc;
      17'd30850: data = 8'h02;
      17'd30851: data = 8'hfe;
      17'd30852: data = 8'h01;
      17'd30853: data = 8'h02;
      17'd30854: data = 8'h02;
      17'd30855: data = 8'h04;
      17'd30856: data = 8'h05;
      17'd30857: data = 8'h05;
      17'd30858: data = 8'h06;
      17'd30859: data = 8'h05;
      17'd30860: data = 8'h01;
      17'd30861: data = 8'h04;
      17'd30862: data = 8'h05;
      17'd30863: data = 8'h01;
      17'd30864: data = 8'h00;
      17'd30865: data = 8'h04;
      17'd30866: data = 8'h04;
      17'd30867: data = 8'h05;
      17'd30868: data = 8'h01;
      17'd30869: data = 8'h02;
      17'd30870: data = 8'h06;
      17'd30871: data = 8'h02;
      17'd30872: data = 8'hfd;
      17'd30873: data = 8'h00;
      17'd30874: data = 8'h09;
      17'd30875: data = 8'h05;
      17'd30876: data = 8'h02;
      17'd30877: data = 8'hfa;
      17'd30878: data = 8'hec;
      17'd30879: data = 8'hfa;
      17'd30880: data = 8'hfe;
      17'd30881: data = 8'h00;
      17'd30882: data = 8'hfe;
      17'd30883: data = 8'he9;
      17'd30884: data = 8'hf5;
      17'd30885: data = 8'h04;
      17'd30886: data = 8'h01;
      17'd30887: data = 8'h06;
      17'd30888: data = 8'h02;
      17'd30889: data = 8'h01;
      17'd30890: data = 8'h05;
      17'd30891: data = 8'h01;
      17'd30892: data = 8'h00;
      17'd30893: data = 8'hef;
      17'd30894: data = 8'hec;
      17'd30895: data = 8'h00;
      17'd30896: data = 8'hfd;
      17'd30897: data = 8'hfc;
      17'd30898: data = 8'h01;
      17'd30899: data = 8'hf2;
      17'd30900: data = 8'hf1;
      17'd30901: data = 8'h01;
      17'd30902: data = 8'hfe;
      17'd30903: data = 8'h01;
      17'd30904: data = 8'h05;
      17'd30905: data = 8'h02;
      17'd30906: data = 8'h01;
      17'd30907: data = 8'hf9;
      17'd30908: data = 8'hf9;
      17'd30909: data = 8'hfa;
      17'd30910: data = 8'hf6;
      17'd30911: data = 8'hfc;
      17'd30912: data = 8'hfa;
      17'd30913: data = 8'hfa;
      17'd30914: data = 8'h02;
      17'd30915: data = 8'h01;
      17'd30916: data = 8'h00;
      17'd30917: data = 8'h02;
      17'd30918: data = 8'h01;
      17'd30919: data = 8'h01;
      17'd30920: data = 8'h02;
      17'd30921: data = 8'h00;
      17'd30922: data = 8'hf9;
      17'd30923: data = 8'hf6;
      17'd30924: data = 8'hf6;
      17'd30925: data = 8'hfd;
      17'd30926: data = 8'hfe;
      17'd30927: data = 8'hf9;
      17'd30928: data = 8'hfc;
      17'd30929: data = 8'hfa;
      17'd30930: data = 8'hfc;
      17'd30931: data = 8'h01;
      17'd30932: data = 8'hfd;
      17'd30933: data = 8'hfa;
      17'd30934: data = 8'hfc;
      17'd30935: data = 8'hfc;
      17'd30936: data = 8'hfd;
      17'd30937: data = 8'hfc;
      17'd30938: data = 8'hfd;
      17'd30939: data = 8'h00;
      17'd30940: data = 8'h00;
      17'd30941: data = 8'h01;
      17'd30942: data = 8'h01;
      17'd30943: data = 8'hfc;
      17'd30944: data = 8'hfd;
      17'd30945: data = 8'hfd;
      17'd30946: data = 8'hf9;
      17'd30947: data = 8'h00;
      17'd30948: data = 8'h05;
      17'd30949: data = 8'h04;
      17'd30950: data = 8'hfd;
      17'd30951: data = 8'hfe;
      17'd30952: data = 8'h0a;
      17'd30953: data = 8'hfe;
      17'd30954: data = 8'hf5;
      17'd30955: data = 8'h00;
      17'd30956: data = 8'h0a;
      17'd30957: data = 8'h05;
      17'd30958: data = 8'h01;
      17'd30959: data = 8'h04;
      17'd30960: data = 8'h01;
      17'd30961: data = 8'h00;
      17'd30962: data = 8'hfe;
      17'd30963: data = 8'h02;
      17'd30964: data = 8'h00;
      17'd30965: data = 8'hf9;
      17'd30966: data = 8'hfa;
      17'd30967: data = 8'hfa;
      17'd30968: data = 8'h00;
      17'd30969: data = 8'hfe;
      17'd30970: data = 8'hf5;
      17'd30971: data = 8'hfc;
      17'd30972: data = 8'h00;
      17'd30973: data = 8'hfc;
      17'd30974: data = 8'hf6;
      17'd30975: data = 8'hfc;
      17'd30976: data = 8'h01;
      17'd30977: data = 8'h01;
      17'd30978: data = 8'hfd;
      17'd30979: data = 8'hfd;
      17'd30980: data = 8'h02;
      17'd30981: data = 8'hfd;
      17'd30982: data = 8'hfa;
      17'd30983: data = 8'hfd;
      17'd30984: data = 8'hfa;
      17'd30985: data = 8'hfa;
      17'd30986: data = 8'hfd;
      17'd30987: data = 8'hfc;
      17'd30988: data = 8'h00;
      17'd30989: data = 8'hfc;
      17'd30990: data = 8'hfd;
      17'd30991: data = 8'h02;
      17'd30992: data = 8'hfc;
      17'd30993: data = 8'hfc;
      17'd30994: data = 8'hf4;
      17'd30995: data = 8'hfe;
      17'd30996: data = 8'h00;
      17'd30997: data = 8'hf5;
      17'd30998: data = 8'h00;
      17'd30999: data = 8'h02;
      17'd31000: data = 8'h06;
      17'd31001: data = 8'h00;
      17'd31002: data = 8'hfd;
      17'd31003: data = 8'hfe;
      17'd31004: data = 8'hfe;
      17'd31005: data = 8'hfd;
      17'd31006: data = 8'hf9;
      17'd31007: data = 8'h00;
      17'd31008: data = 8'h00;
      17'd31009: data = 8'h00;
      17'd31010: data = 8'h0a;
      17'd31011: data = 8'h02;
      17'd31012: data = 8'h00;
      17'd31013: data = 8'h01;
      17'd31014: data = 8'h05;
      17'd31015: data = 8'h0c;
      17'd31016: data = 8'h01;
      17'd31017: data = 8'hfc;
      17'd31018: data = 8'hfc;
      17'd31019: data = 8'h06;
      17'd31020: data = 8'h04;
      17'd31021: data = 8'h00;
      17'd31022: data = 8'h02;
      17'd31023: data = 8'h04;
      17'd31024: data = 8'h05;
      17'd31025: data = 8'hf9;
      17'd31026: data = 8'h00;
      17'd31027: data = 8'h0a;
      17'd31028: data = 8'h00;
      17'd31029: data = 8'h05;
      17'd31030: data = 8'hfe;
      17'd31031: data = 8'hfe;
      17'd31032: data = 8'h02;
      17'd31033: data = 8'hf6;
      17'd31034: data = 8'hfa;
      17'd31035: data = 8'hfe;
      17'd31036: data = 8'hf6;
      17'd31037: data = 8'hf9;
      17'd31038: data = 8'hf5;
      17'd31039: data = 8'hfd;
      17'd31040: data = 8'h00;
      17'd31041: data = 8'hf6;
      17'd31042: data = 8'h05;
      17'd31043: data = 8'h0a;
      17'd31044: data = 8'h05;
      17'd31045: data = 8'h02;
      17'd31046: data = 8'hf9;
      17'd31047: data = 8'hfd;
      17'd31048: data = 8'hfe;
      17'd31049: data = 8'hf5;
      17'd31050: data = 8'hfa;
      17'd31051: data = 8'hf9;
      17'd31052: data = 8'hfa;
      17'd31053: data = 8'h02;
      17'd31054: data = 8'hfa;
      17'd31055: data = 8'hfc;
      17'd31056: data = 8'h05;
      17'd31057: data = 8'h04;
      17'd31058: data = 8'h01;
      17'd31059: data = 8'h01;
      17'd31060: data = 8'h06;
      17'd31061: data = 8'h05;
      17'd31062: data = 8'hfe;
      17'd31063: data = 8'h0c;
      17'd31064: data = 8'h0c;
      17'd31065: data = 8'h00;
      17'd31066: data = 8'h06;
      17'd31067: data = 8'hfe;
      17'd31068: data = 8'hfc;
      17'd31069: data = 8'h00;
      17'd31070: data = 8'hfa;
      17'd31071: data = 8'h05;
      17'd31072: data = 8'h02;
      17'd31073: data = 8'hfc;
      17'd31074: data = 8'h02;
      17'd31075: data = 8'h00;
      17'd31076: data = 8'h05;
      17'd31077: data = 8'h05;
      17'd31078: data = 8'h01;
      17'd31079: data = 8'h11;
      17'd31080: data = 8'h02;
      17'd31081: data = 8'hfe;
      17'd31082: data = 8'h06;
      17'd31083: data = 8'h00;
      17'd31084: data = 8'hfc;
      17'd31085: data = 8'hfe;
      17'd31086: data = 8'hf2;
      17'd31087: data = 8'hfa;
      17'd31088: data = 8'hfd;
      17'd31089: data = 8'hfe;
      17'd31090: data = 8'h0a;
      17'd31091: data = 8'h04;
      17'd31092: data = 8'h0a;
      17'd31093: data = 8'h0c;
      17'd31094: data = 8'hf6;
      17'd31095: data = 8'hfc;
      17'd31096: data = 8'hfd;
      17'd31097: data = 8'hf5;
      17'd31098: data = 8'h05;
      17'd31099: data = 8'h01;
      17'd31100: data = 8'h06;
      17'd31101: data = 8'h11;
      17'd31102: data = 8'h04;
      17'd31103: data = 8'h02;
      17'd31104: data = 8'h00;
      17'd31105: data = 8'h00;
      17'd31106: data = 8'hf2;
      17'd31107: data = 8'hf1;
      17'd31108: data = 8'hfe;
      17'd31109: data = 8'hfd;
      17'd31110: data = 8'hf6;
      17'd31111: data = 8'h00;
      17'd31112: data = 8'h02;
      17'd31113: data = 8'hfd;
      17'd31114: data = 8'h04;
      17'd31115: data = 8'h01;
      17'd31116: data = 8'h05;
      17'd31117: data = 8'h04;
      17'd31118: data = 8'hf6;
      17'd31119: data = 8'hfe;
      17'd31120: data = 8'hf9;
      17'd31121: data = 8'hfd;
      17'd31122: data = 8'h00;
      17'd31123: data = 8'hf2;
      17'd31124: data = 8'h02;
      17'd31125: data = 8'h05;
      17'd31126: data = 8'hfd;
      17'd31127: data = 8'h09;
      17'd31128: data = 8'h04;
      17'd31129: data = 8'h05;
      17'd31130: data = 8'h0c;
      17'd31131: data = 8'hfc;
      17'd31132: data = 8'hfd;
      17'd31133: data = 8'hfd;
      17'd31134: data = 8'hf2;
      17'd31135: data = 8'hfa;
      17'd31136: data = 8'hf2;
      17'd31137: data = 8'hf2;
      17'd31138: data = 8'h02;
      17'd31139: data = 8'hfc;
      17'd31140: data = 8'h01;
      17'd31141: data = 8'h0d;
      17'd31142: data = 8'hfe;
      17'd31143: data = 8'h04;
      17'd31144: data = 8'h09;
      17'd31145: data = 8'hfe;
      17'd31146: data = 8'h00;
      17'd31147: data = 8'hf5;
      17'd31148: data = 8'hfe;
      17'd31149: data = 8'h05;
      17'd31150: data = 8'hfd;
      17'd31151: data = 8'h05;
      17'd31152: data = 8'hf4;
      17'd31153: data = 8'hf6;
      17'd31154: data = 8'h04;
      17'd31155: data = 8'h01;
      17'd31156: data = 8'hfc;
      17'd31157: data = 8'hf9;
      17'd31158: data = 8'h05;
      17'd31159: data = 8'h05;
      17'd31160: data = 8'h09;
      17'd31161: data = 8'h0d;
      17'd31162: data = 8'h09;
      17'd31163: data = 8'h09;
      17'd31164: data = 8'h00;
      17'd31165: data = 8'hfc;
      17'd31166: data = 8'hf5;
      17'd31167: data = 8'hf4;
      17'd31168: data = 8'hfc;
      17'd31169: data = 8'h01;
      17'd31170: data = 8'hfc;
      17'd31171: data = 8'hf6;
      17'd31172: data = 8'hf9;
      17'd31173: data = 8'hfd;
      17'd31174: data = 8'hfc;
      17'd31175: data = 8'h01;
      17'd31176: data = 8'hfe;
      17'd31177: data = 8'hfe;
      17'd31178: data = 8'h09;
      17'd31179: data = 8'h0a;
      17'd31180: data = 8'h09;
      17'd31181: data = 8'h04;
      17'd31182: data = 8'h0c;
      17'd31183: data = 8'hfe;
      17'd31184: data = 8'h00;
      17'd31185: data = 8'hfe;
      17'd31186: data = 8'hed;
      17'd31187: data = 8'hf6;
      17'd31188: data = 8'hfe;
      17'd31189: data = 8'hf6;
      17'd31190: data = 8'hfa;
      17'd31191: data = 8'h01;
      17'd31192: data = 8'h05;
      17'd31193: data = 8'h09;
      17'd31194: data = 8'h01;
      17'd31195: data = 8'hfd;
      17'd31196: data = 8'hfa;
      17'd31197: data = 8'hf5;
      17'd31198: data = 8'hfd;
      17'd31199: data = 8'hf9;
      17'd31200: data = 8'h01;
      17'd31201: data = 8'hfe;
      17'd31202: data = 8'hf9;
      17'd31203: data = 8'h02;
      17'd31204: data = 8'h00;
      17'd31205: data = 8'h02;
      17'd31206: data = 8'hfc;
      17'd31207: data = 8'hf5;
      17'd31208: data = 8'h02;
      17'd31209: data = 8'hfe;
      17'd31210: data = 8'hf4;
      17'd31211: data = 8'h04;
      17'd31212: data = 8'h04;
      17'd31213: data = 8'hfd;
      17'd31214: data = 8'h0d;
      17'd31215: data = 8'h02;
      17'd31216: data = 8'hf9;
      17'd31217: data = 8'h0e;
      17'd31218: data = 8'h05;
      17'd31219: data = 8'hfd;
      17'd31220: data = 8'h0a;
      17'd31221: data = 8'h05;
      17'd31222: data = 8'h01;
      17'd31223: data = 8'h0a;
      17'd31224: data = 8'h0a;
      17'd31225: data = 8'h00;
      17'd31226: data = 8'hfc;
      17'd31227: data = 8'hf9;
      17'd31228: data = 8'hf9;
      17'd31229: data = 8'heb;
      17'd31230: data = 8'hf6;
      17'd31231: data = 8'h04;
      17'd31232: data = 8'hed;
      17'd31233: data = 8'hfd;
      17'd31234: data = 8'h0a;
      17'd31235: data = 8'h01;
      17'd31236: data = 8'hfd;
      17'd31237: data = 8'h00;
      17'd31238: data = 8'h04;
      17'd31239: data = 8'hf4;
      17'd31240: data = 8'h02;
      17'd31241: data = 8'h0a;
      17'd31242: data = 8'hf2;
      17'd31243: data = 8'hfe;
      17'd31244: data = 8'h06;
      17'd31245: data = 8'h01;
      17'd31246: data = 8'h00;
      17'd31247: data = 8'h02;
      17'd31248: data = 8'h05;
      17'd31249: data = 8'h00;
      17'd31250: data = 8'h04;
      17'd31251: data = 8'hf9;
      17'd31252: data = 8'hf1;
      17'd31253: data = 8'hfe;
      17'd31254: data = 8'h01;
      17'd31255: data = 8'hfa;
      17'd31256: data = 8'hfa;
      17'd31257: data = 8'hfc;
      17'd31258: data = 8'hf5;
      17'd31259: data = 8'h00;
      17'd31260: data = 8'h01;
      17'd31261: data = 8'h02;
      17'd31262: data = 8'h0d;
      17'd31263: data = 8'h05;
      17'd31264: data = 8'h04;
      17'd31265: data = 8'h02;
      17'd31266: data = 8'h05;
      17'd31267: data = 8'h06;
      17'd31268: data = 8'h01;
      17'd31269: data = 8'h0a;
      17'd31270: data = 8'h06;
      17'd31271: data = 8'h05;
      17'd31272: data = 8'h02;
      17'd31273: data = 8'h01;
      17'd31274: data = 8'h02;
      17'd31275: data = 8'hfc;
      17'd31276: data = 8'hfc;
      17'd31277: data = 8'h06;
      17'd31278: data = 8'hfd;
      17'd31279: data = 8'hfe;
      17'd31280: data = 8'hfd;
      17'd31281: data = 8'hf5;
      17'd31282: data = 8'h06;
      17'd31283: data = 8'hfc;
      17'd31284: data = 8'hf5;
      17'd31285: data = 8'h02;
      17'd31286: data = 8'hfc;
      17'd31287: data = 8'h04;
      17'd31288: data = 8'h00;
      17'd31289: data = 8'he5;
      17'd31290: data = 8'h00;
      17'd31291: data = 8'h02;
      17'd31292: data = 8'hf9;
      17'd31293: data = 8'h0a;
      17'd31294: data = 8'h00;
      17'd31295: data = 8'hfc;
      17'd31296: data = 8'h00;
      17'd31297: data = 8'hfd;
      17'd31298: data = 8'h13;
      17'd31299: data = 8'h0d;
      17'd31300: data = 8'hfe;
      17'd31301: data = 8'h0a;
      17'd31302: data = 8'h0e;
      17'd31303: data = 8'h09;
      17'd31304: data = 8'h02;
      17'd31305: data = 8'hfe;
      17'd31306: data = 8'hfd;
      17'd31307: data = 8'hfd;
      17'd31308: data = 8'he9;
      17'd31309: data = 8'hf1;
      17'd31310: data = 8'hfd;
      17'd31311: data = 8'hf6;
      17'd31312: data = 8'h09;
      17'd31313: data = 8'h04;
      17'd31314: data = 8'h05;
      17'd31315: data = 8'h12;
      17'd31316: data = 8'h15;
      17'd31317: data = 8'h0e;
      17'd31318: data = 8'h00;
      17'd31319: data = 8'h05;
      17'd31320: data = 8'h0a;
      17'd31321: data = 8'h01;
      17'd31322: data = 8'hf9;
      17'd31323: data = 8'hf4;
      17'd31324: data = 8'h01;
      17'd31325: data = 8'hf4;
      17'd31326: data = 8'hf9;
      17'd31327: data = 8'h0d;
      17'd31328: data = 8'hf1;
      17'd31329: data = 8'h06;
      17'd31330: data = 8'h19;
      17'd31331: data = 8'hfc;
      17'd31332: data = 8'h0a;
      17'd31333: data = 8'hfc;
      17'd31334: data = 8'heb;
      17'd31335: data = 8'hf9;
      17'd31336: data = 8'hf9;
      17'd31337: data = 8'h0a;
      17'd31338: data = 8'h05;
      17'd31339: data = 8'hfc;
      17'd31340: data = 8'h0c;
      17'd31341: data = 8'hfa;
      17'd31342: data = 8'hf9;
      17'd31343: data = 8'h0a;
      17'd31344: data = 8'hf2;
      17'd31345: data = 8'hfc;
      17'd31346: data = 8'h00;
      17'd31347: data = 8'hf1;
      17'd31348: data = 8'hfa;
      17'd31349: data = 8'hf4;
      17'd31350: data = 8'h00;
      17'd31351: data = 8'h02;
      17'd31352: data = 8'hf9;
      17'd31353: data = 8'h01;
      17'd31354: data = 8'hfa;
      17'd31355: data = 8'hf6;
      17'd31356: data = 8'h05;
      17'd31357: data = 8'h0d;
      17'd31358: data = 8'h0c;
      17'd31359: data = 8'h05;
      17'd31360: data = 8'h0d;
      17'd31361: data = 8'h04;
      17'd31362: data = 8'heb;
      17'd31363: data = 8'hec;
      17'd31364: data = 8'hf6;
      17'd31365: data = 8'hf1;
      17'd31366: data = 8'hf5;
      17'd31367: data = 8'hfd;
      17'd31368: data = 8'hfd;
      17'd31369: data = 8'h0a;
      17'd31370: data = 8'h0c;
      17'd31371: data = 8'hfe;
      17'd31372: data = 8'h05;
      17'd31373: data = 8'h02;
      17'd31374: data = 8'h01;
      17'd31375: data = 8'h02;
      17'd31376: data = 8'hfa;
      17'd31377: data = 8'hfd;
      17'd31378: data = 8'hf9;
      17'd31379: data = 8'h00;
      17'd31380: data = 8'hfc;
      17'd31381: data = 8'hfa;
      17'd31382: data = 8'h01;
      17'd31383: data = 8'hfc;
      17'd31384: data = 8'hfc;
      17'd31385: data = 8'h02;
      17'd31386: data = 8'hfc;
      17'd31387: data = 8'hf2;
      17'd31388: data = 8'h02;
      17'd31389: data = 8'hf9;
      17'd31390: data = 8'h09;
      17'd31391: data = 8'h06;
      17'd31392: data = 8'hf5;
      17'd31393: data = 8'h0d;
      17'd31394: data = 8'hf6;
      17'd31395: data = 8'h02;
      17'd31396: data = 8'h0c;
      17'd31397: data = 8'he5;
      17'd31398: data = 8'hfd;
      17'd31399: data = 8'h00;
      17'd31400: data = 8'hf4;
      17'd31401: data = 8'h06;
      17'd31402: data = 8'hed;
      17'd31403: data = 8'hf5;
      17'd31404: data = 8'h00;
      17'd31405: data = 8'hef;
      17'd31406: data = 8'h00;
      17'd31407: data = 8'hfc;
      17'd31408: data = 8'h00;
      17'd31409: data = 8'h09;
      17'd31410: data = 8'hf6;
      17'd31411: data = 8'h0e;
      17'd31412: data = 8'h0e;
      17'd31413: data = 8'hfa;
      17'd31414: data = 8'h06;
      17'd31415: data = 8'hfd;
      17'd31416: data = 8'h01;
      17'd31417: data = 8'h05;
      17'd31418: data = 8'he3;
      17'd31419: data = 8'hf5;
      17'd31420: data = 8'h04;
      17'd31421: data = 8'hf2;
      17'd31422: data = 8'hfc;
      17'd31423: data = 8'hfe;
      17'd31424: data = 8'h01;
      17'd31425: data = 8'h01;
      17'd31426: data = 8'hfe;
      17'd31427: data = 8'h0c;
      17'd31428: data = 8'hfd;
      17'd31429: data = 8'hf5;
      17'd31430: data = 8'h05;
      17'd31431: data = 8'hfd;
      17'd31432: data = 8'hfd;
      17'd31433: data = 8'hf6;
      17'd31434: data = 8'hf5;
      17'd31435: data = 8'h04;
      17'd31436: data = 8'hfd;
      17'd31437: data = 8'hfe;
      17'd31438: data = 8'h05;
      17'd31439: data = 8'h00;
      17'd31440: data = 8'h11;
      17'd31441: data = 8'h06;
      17'd31442: data = 8'hf5;
      17'd31443: data = 8'hfa;
      17'd31444: data = 8'hf1;
      17'd31445: data = 8'hf9;
      17'd31446: data = 8'hf9;
      17'd31447: data = 8'hf1;
      17'd31448: data = 8'h00;
      17'd31449: data = 8'hfe;
      17'd31450: data = 8'hfe;
      17'd31451: data = 8'h0c;
      17'd31452: data = 8'h00;
      17'd31453: data = 8'hfe;
      17'd31454: data = 8'h0d;
      17'd31455: data = 8'h02;
      17'd31456: data = 8'h0d;
      17'd31457: data = 8'h0a;
      17'd31458: data = 8'hfa;
      17'd31459: data = 8'hfe;
      17'd31460: data = 8'hf9;
      17'd31461: data = 8'hfe;
      17'd31462: data = 8'hf4;
      17'd31463: data = 8'hfa;
      17'd31464: data = 8'h09;
      17'd31465: data = 8'hf9;
      17'd31466: data = 8'h04;
      17'd31467: data = 8'h12;
      17'd31468: data = 8'h01;
      17'd31469: data = 8'h01;
      17'd31470: data = 8'h09;
      17'd31471: data = 8'h01;
      17'd31472: data = 8'hfe;
      17'd31473: data = 8'hfc;
      17'd31474: data = 8'h00;
      17'd31475: data = 8'hfc;
      17'd31476: data = 8'hf2;
      17'd31477: data = 8'hfa;
      17'd31478: data = 8'hf1;
      17'd31479: data = 8'hfa;
      17'd31480: data = 8'hfd;
      17'd31481: data = 8'hf2;
      17'd31482: data = 8'hfd;
      17'd31483: data = 8'h00;
      17'd31484: data = 8'h0a;
      17'd31485: data = 8'h13;
      17'd31486: data = 8'h02;
      17'd31487: data = 8'h05;
      17'd31488: data = 8'h0a;
      17'd31489: data = 8'hfe;
      17'd31490: data = 8'h01;
      17'd31491: data = 8'hf4;
      17'd31492: data = 8'hed;
      17'd31493: data = 8'h01;
      17'd31494: data = 8'hfa;
      17'd31495: data = 8'hfe;
      17'd31496: data = 8'h09;
      17'd31497: data = 8'hfa;
      17'd31498: data = 8'hfd;
      17'd31499: data = 8'h06;
      17'd31500: data = 8'h05;
      17'd31501: data = 8'h02;
      17'd31502: data = 8'hfe;
      17'd31503: data = 8'hf9;
      17'd31504: data = 8'hfc;
      17'd31505: data = 8'hf9;
      17'd31506: data = 8'h01;
      17'd31507: data = 8'hfe;
      17'd31508: data = 8'hfc;
      17'd31509: data = 8'h0e;
      17'd31510: data = 8'h02;
      17'd31511: data = 8'hfa;
      17'd31512: data = 8'h00;
      17'd31513: data = 8'h01;
      17'd31514: data = 8'h02;
      17'd31515: data = 8'hfe;
      17'd31516: data = 8'hfd;
      17'd31517: data = 8'hfa;
      17'd31518: data = 8'hf5;
      17'd31519: data = 8'hfa;
      17'd31520: data = 8'h00;
      17'd31521: data = 8'hfe;
      17'd31522: data = 8'h06;
      17'd31523: data = 8'h0e;
      17'd31524: data = 8'h0c;
      17'd31525: data = 8'h0d;
      17'd31526: data = 8'h05;
      17'd31527: data = 8'h02;
      17'd31528: data = 8'hfd;
      17'd31529: data = 8'hfd;
      17'd31530: data = 8'hf1;
      17'd31531: data = 8'he4;
      17'd31532: data = 8'hef;
      17'd31533: data = 8'hf6;
      17'd31534: data = 8'hf1;
      17'd31535: data = 8'hfa;
      17'd31536: data = 8'h0a;
      17'd31537: data = 8'h06;
      17'd31538: data = 8'h16;
      17'd31539: data = 8'h1f;
      17'd31540: data = 8'h12;
      17'd31541: data = 8'h04;
      17'd31542: data = 8'h00;
      17'd31543: data = 8'h09;
      17'd31544: data = 8'hf2;
      17'd31545: data = 8'hed;
      17'd31546: data = 8'hf6;
      17'd31547: data = 8'hec;
      17'd31548: data = 8'h00;
      17'd31549: data = 8'h06;
      17'd31550: data = 8'hf6;
      17'd31551: data = 8'hfd;
      17'd31552: data = 8'h0e;
      17'd31553: data = 8'h15;
      17'd31554: data = 8'h15;
      17'd31555: data = 8'h0c;
      17'd31556: data = 8'h01;
      17'd31557: data = 8'hfc;
      17'd31558: data = 8'hf6;
      17'd31559: data = 8'hfc;
      17'd31560: data = 8'hf6;
      17'd31561: data = 8'hf6;
      17'd31562: data = 8'hfe;
      17'd31563: data = 8'h02;
      17'd31564: data = 8'h04;
      17'd31565: data = 8'h05;
      17'd31566: data = 8'h0c;
      17'd31567: data = 8'h0d;
      17'd31568: data = 8'h06;
      17'd31569: data = 8'h04;
      17'd31570: data = 8'h00;
      17'd31571: data = 8'hf5;
      17'd31572: data = 8'hf5;
      17'd31573: data = 8'hfc;
      17'd31574: data = 8'h06;
      17'd31575: data = 8'h0a;
      17'd31576: data = 8'h00;
      17'd31577: data = 8'hfa;
      17'd31578: data = 8'h02;
      17'd31579: data = 8'h01;
      17'd31580: data = 8'hfa;
      17'd31581: data = 8'h01;
      17'd31582: data = 8'h01;
      17'd31583: data = 8'h04;
      17'd31584: data = 8'h02;
      17'd31585: data = 8'hf4;
      17'd31586: data = 8'hf9;
      17'd31587: data = 8'hf5;
      17'd31588: data = 8'h01;
      17'd31589: data = 8'h0d;
      17'd31590: data = 8'hfd;
      17'd31591: data = 8'h01;
      17'd31592: data = 8'h04;
      17'd31593: data = 8'hf9;
      17'd31594: data = 8'hfd;
      17'd31595: data = 8'h04;
      17'd31596: data = 8'hfa;
      17'd31597: data = 8'hf6;
      17'd31598: data = 8'hfc;
      17'd31599: data = 8'hfc;
      17'd31600: data = 8'hfc;
      17'd31601: data = 8'hfc;
      17'd31602: data = 8'h00;
      17'd31603: data = 8'h05;
      17'd31604: data = 8'h06;
      17'd31605: data = 8'h0d;
      17'd31606: data = 8'h09;
      17'd31607: data = 8'hfa;
      17'd31608: data = 8'h00;
      17'd31609: data = 8'hfd;
      17'd31610: data = 8'hf9;
      17'd31611: data = 8'h00;
      17'd31612: data = 8'hfd;
      17'd31613: data = 8'hf6;
      17'd31614: data = 8'hfc;
      17'd31615: data = 8'h09;
      17'd31616: data = 8'h04;
      17'd31617: data = 8'h00;
      17'd31618: data = 8'h09;
      17'd31619: data = 8'h0a;
      17'd31620: data = 8'h06;
      17'd31621: data = 8'h01;
      17'd31622: data = 8'h01;
      17'd31623: data = 8'h00;
      17'd31624: data = 8'hf6;
      17'd31625: data = 8'hf1;
      17'd31626: data = 8'hef;
      17'd31627: data = 8'hf9;
      17'd31628: data = 8'h01;
      17'd31629: data = 8'hf5;
      17'd31630: data = 8'hf9;
      17'd31631: data = 8'hfe;
      17'd31632: data = 8'hfd;
      17'd31633: data = 8'hfe;
      17'd31634: data = 8'h06;
      17'd31635: data = 8'h11;
      17'd31636: data = 8'h09;
      17'd31637: data = 8'h00;
      17'd31638: data = 8'hfa;
      17'd31639: data = 8'hf9;
      17'd31640: data = 8'hf2;
      17'd31641: data = 8'hf1;
      17'd31642: data = 8'hf2;
      17'd31643: data = 8'hf4;
      17'd31644: data = 8'hfe;
      17'd31645: data = 8'h06;
      17'd31646: data = 8'h05;
      17'd31647: data = 8'h0c;
      17'd31648: data = 8'h0a;
      17'd31649: data = 8'h0c;
      17'd31650: data = 8'h0e;
      17'd31651: data = 8'h06;
      17'd31652: data = 8'h01;
      17'd31653: data = 8'hf6;
      17'd31654: data = 8'hed;
      17'd31655: data = 8'hf2;
      17'd31656: data = 8'hf9;
      17'd31657: data = 8'hfd;
      17'd31658: data = 8'h00;
      17'd31659: data = 8'hfc;
      17'd31660: data = 8'h01;
      17'd31661: data = 8'h06;
      17'd31662: data = 8'h05;
      17'd31663: data = 8'h06;
      17'd31664: data = 8'h05;
      17'd31665: data = 8'h05;
      17'd31666: data = 8'h05;
      17'd31667: data = 8'hfe;
      17'd31668: data = 8'hfe;
      17'd31669: data = 8'hfd;
      17'd31670: data = 8'hf4;
      17'd31671: data = 8'hf9;
      17'd31672: data = 8'hfa;
      17'd31673: data = 8'hf9;
      17'd31674: data = 8'hfe;
      17'd31675: data = 8'hfd;
      17'd31676: data = 8'hfe;
      17'd31677: data = 8'hfe;
      17'd31678: data = 8'hfa;
      17'd31679: data = 8'h00;
      17'd31680: data = 8'hfa;
      17'd31681: data = 8'hf2;
      17'd31682: data = 8'hf9;
      17'd31683: data = 8'hf6;
      17'd31684: data = 8'hf6;
      17'd31685: data = 8'hf9;
      17'd31686: data = 8'hfd;
      17'd31687: data = 8'h04;
      17'd31688: data = 8'h06;
      17'd31689: data = 8'h06;
      17'd31690: data = 8'h05;
      17'd31691: data = 8'h05;
      17'd31692: data = 8'hfc;
      17'd31693: data = 8'hf5;
      17'd31694: data = 8'hfc;
      17'd31695: data = 8'hf6;
      17'd31696: data = 8'hf2;
      17'd31697: data = 8'hfa;
      17'd31698: data = 8'hf9;
      17'd31699: data = 8'hfa;
      17'd31700: data = 8'h04;
      17'd31701: data = 8'h0a;
      17'd31702: data = 8'h09;
      17'd31703: data = 8'h0c;
      17'd31704: data = 8'h12;
      17'd31705: data = 8'h0c;
      17'd31706: data = 8'h04;
      17'd31707: data = 8'h02;
      17'd31708: data = 8'hfc;
      17'd31709: data = 8'hf4;
      17'd31710: data = 8'hf4;
      17'd31711: data = 8'hf5;
      17'd31712: data = 8'hf4;
      17'd31713: data = 8'hf5;
      17'd31714: data = 8'hfa;
      17'd31715: data = 8'hfe;
      17'd31716: data = 8'h01;
      17'd31717: data = 8'h05;
      17'd31718: data = 8'h05;
      17'd31719: data = 8'hfd;
      17'd31720: data = 8'h00;
      17'd31721: data = 8'h01;
      17'd31722: data = 8'hfe;
      17'd31723: data = 8'h01;
      17'd31724: data = 8'hfd;
      17'd31725: data = 8'hfc;
      17'd31726: data = 8'h00;
      17'd31727: data = 8'h04;
      17'd31728: data = 8'h09;
      17'd31729: data = 8'h02;
      17'd31730: data = 8'hfe;
      17'd31731: data = 8'h00;
      17'd31732: data = 8'hfa;
      17'd31733: data = 8'hfd;
      17'd31734: data = 8'hfd;
      17'd31735: data = 8'hfd;
      17'd31736: data = 8'hfd;
      17'd31737: data = 8'hf6;
      17'd31738: data = 8'hfe;
      17'd31739: data = 8'hfe;
      17'd31740: data = 8'hfd;
      17'd31741: data = 8'h05;
      17'd31742: data = 8'h05;
      17'd31743: data = 8'h06;
      17'd31744: data = 8'h0a;
      17'd31745: data = 8'h04;
      17'd31746: data = 8'h02;
      17'd31747: data = 8'hfc;
      17'd31748: data = 8'hf9;
      17'd31749: data = 8'hfd;
      17'd31750: data = 8'hfe;
      17'd31751: data = 8'hfd;
      17'd31752: data = 8'hfa;
      17'd31753: data = 8'hf9;
      17'd31754: data = 8'hf9;
      17'd31755: data = 8'hfe;
      17'd31756: data = 8'h04;
      17'd31757: data = 8'h06;
      17'd31758: data = 8'h09;
      17'd31759: data = 8'h05;
      17'd31760: data = 8'h02;
      17'd31761: data = 8'h01;
      17'd31762: data = 8'h02;
      17'd31763: data = 8'h00;
      17'd31764: data = 8'hfa;
      17'd31765: data = 8'hfa;
      17'd31766: data = 8'h00;
      17'd31767: data = 8'h01;
      17'd31768: data = 8'h00;
      17'd31769: data = 8'h01;
      17'd31770: data = 8'h02;
      17'd31771: data = 8'h02;
      17'd31772: data = 8'h04;
      17'd31773: data = 8'h09;
      17'd31774: data = 8'h06;
      17'd31775: data = 8'hfe;
      17'd31776: data = 8'hfa;
      17'd31777: data = 8'hfd;
      17'd31778: data = 8'hfd;
      17'd31779: data = 8'h01;
      17'd31780: data = 8'hfe;
      17'd31781: data = 8'h00;
      17'd31782: data = 8'h04;
      17'd31783: data = 8'h01;
      17'd31784: data = 8'h02;
      17'd31785: data = 8'h01;
      17'd31786: data = 8'h04;
      17'd31787: data = 8'h01;
      17'd31788: data = 8'hfc;
      17'd31789: data = 8'hfe;
      17'd31790: data = 8'hfe;
      17'd31791: data = 8'hfe;
      17'd31792: data = 8'hfa;
      17'd31793: data = 8'hf9;
      17'd31794: data = 8'hfc;
      17'd31795: data = 8'h00;
      17'd31796: data = 8'h02;
      17'd31797: data = 8'h01;
      17'd31798: data = 8'h04;
      17'd31799: data = 8'h04;
      17'd31800: data = 8'h01;
      17'd31801: data = 8'hfe;
      17'd31802: data = 8'hfe;
      17'd31803: data = 8'hfe;
      17'd31804: data = 8'hfe;
      17'd31805: data = 8'hf9;
      17'd31806: data = 8'hf9;
      17'd31807: data = 8'hf9;
      17'd31808: data = 8'hf9;
      17'd31809: data = 8'hfd;
      17'd31810: data = 8'hfc;
      17'd31811: data = 8'h02;
      17'd31812: data = 8'h04;
      17'd31813: data = 8'h01;
      17'd31814: data = 8'hfe;
      17'd31815: data = 8'hfe;
      17'd31816: data = 8'h02;
      17'd31817: data = 8'hfd;
      17'd31818: data = 8'hfc;
      17'd31819: data = 8'hfd;
      17'd31820: data = 8'h02;
      17'd31821: data = 8'h00;
      17'd31822: data = 8'hf9;
      17'd31823: data = 8'h00;
      17'd31824: data = 8'h01;
      17'd31825: data = 8'hfc;
      17'd31826: data = 8'hfe;
      17'd31827: data = 8'h02;
      17'd31828: data = 8'h05;
      17'd31829: data = 8'h05;
      17'd31830: data = 8'h05;
      17'd31831: data = 8'h09;
      17'd31832: data = 8'h04;
      17'd31833: data = 8'h05;
      17'd31834: data = 8'h05;
      17'd31835: data = 8'hfe;
      17'd31836: data = 8'hfc;
      17'd31837: data = 8'hfc;
      17'd31838: data = 8'hfe;
      17'd31839: data = 8'hfc;
      17'd31840: data = 8'hfe;
      17'd31841: data = 8'hfd;
      17'd31842: data = 8'hfe;
      17'd31843: data = 8'hfc;
      17'd31844: data = 8'h01;
      17'd31845: data = 8'h05;
      17'd31846: data = 8'hfd;
      17'd31847: data = 8'h00;
      17'd31848: data = 8'h01;
      17'd31849: data = 8'h02;
      17'd31850: data = 8'h01;
      17'd31851: data = 8'h00;
      17'd31852: data = 8'hfd;
      17'd31853: data = 8'hfc;
      17'd31854: data = 8'hfa;
      17'd31855: data = 8'hf6;
      17'd31856: data = 8'hf6;
      17'd31857: data = 8'hf5;
      17'd31858: data = 8'hfa;
      17'd31859: data = 8'hf6;
      17'd31860: data = 8'hfa;
      17'd31861: data = 8'h01;
      17'd31862: data = 8'h00;
      17'd31863: data = 8'hfe;
      17'd31864: data = 8'h04;
      17'd31865: data = 8'h02;
      17'd31866: data = 8'h01;
      17'd31867: data = 8'h02;
      17'd31868: data = 8'h04;
      17'd31869: data = 8'h00;
      17'd31870: data = 8'hfe;
      17'd31871: data = 8'h05;
      17'd31872: data = 8'h01;
      17'd31873: data = 8'h00;
      17'd31874: data = 8'h05;
      17'd31875: data = 8'h06;
      17'd31876: data = 8'h04;
      17'd31877: data = 8'hfe;
      17'd31878: data = 8'hfc;
      17'd31879: data = 8'hf5;
      17'd31880: data = 8'he7;
      17'd31881: data = 8'he0;
      17'd31882: data = 8'he4;
      17'd31883: data = 8'he7;
      17'd31884: data = 8'hed;
      17'd31885: data = 8'hf2;
      17'd31886: data = 8'h04;
      17'd31887: data = 8'h11;
      17'd31888: data = 8'h13;
      17'd31889: data = 8'h1e;
      17'd31890: data = 8'h1f;
      17'd31891: data = 8'h1f;
      17'd31892: data = 8'h1e;
      17'd31893: data = 8'h1a;
      17'd31894: data = 8'h12;
      17'd31895: data = 8'h0c;
      17'd31896: data = 8'h05;
      17'd31897: data = 8'hfe;
      17'd31898: data = 8'hfc;
      17'd31899: data = 8'hfd;
      17'd31900: data = 8'hfe;
      17'd31901: data = 8'hf5;
      17'd31902: data = 8'hf9;
      17'd31903: data = 8'h02;
      17'd31904: data = 8'hfa;
      17'd31905: data = 8'hf5;
      17'd31906: data = 8'hfa;
      17'd31907: data = 8'hf9;
      17'd31908: data = 8'hf4;
      17'd31909: data = 8'hef;
      17'd31910: data = 8'hf4;
      17'd31911: data = 8'hf6;
      17'd31912: data = 8'hf6;
      17'd31913: data = 8'hfc;
      17'd31914: data = 8'hf9;
      17'd31915: data = 8'hfd;
      17'd31916: data = 8'hfd;
      17'd31917: data = 8'hf1;
      17'd31918: data = 8'heb;
      17'd31919: data = 8'hef;
      17'd31920: data = 8'hf1;
      17'd31921: data = 8'he4;
      17'd31922: data = 8'he7;
      17'd31923: data = 8'hf9;
      17'd31924: data = 8'hf6;
      17'd31925: data = 8'hf4;
      17'd31926: data = 8'hfe;
      17'd31927: data = 8'h04;
      17'd31928: data = 8'h02;
      17'd31929: data = 8'h01;
      17'd31930: data = 8'h05;
      17'd31931: data = 8'h09;
      17'd31932: data = 8'h05;
      17'd31933: data = 8'h02;
      17'd31934: data = 8'h01;
      17'd31935: data = 8'h04;
      17'd31936: data = 8'h09;
      17'd31937: data = 8'h04;
      17'd31938: data = 8'h02;
      17'd31939: data = 8'h09;
      17'd31940: data = 8'h0c;
      17'd31941: data = 8'h05;
      17'd31942: data = 8'h01;
      17'd31943: data = 8'h09;
      17'd31944: data = 8'h06;
      17'd31945: data = 8'h02;
      17'd31946: data = 8'h09;
      17'd31947: data = 8'h11;
      17'd31948: data = 8'h12;
      17'd31949: data = 8'h0d;
      17'd31950: data = 8'h11;
      17'd31951: data = 8'h16;
      17'd31952: data = 8'h11;
      17'd31953: data = 8'h0a;
      17'd31954: data = 8'h0c;
      17'd31955: data = 8'h0a;
      17'd31956: data = 8'h0a;
      17'd31957: data = 8'h06;
      17'd31958: data = 8'h04;
      17'd31959: data = 8'h05;
      17'd31960: data = 8'h05;
      17'd31961: data = 8'h06;
      17'd31962: data = 8'h02;
      17'd31963: data = 8'h02;
      17'd31964: data = 8'h04;
      17'd31965: data = 8'h00;
      17'd31966: data = 8'hfd;
      17'd31967: data = 8'hfd;
      17'd31968: data = 8'h00;
      17'd31969: data = 8'hfc;
      17'd31970: data = 8'hf6;
      17'd31971: data = 8'hfe;
      17'd31972: data = 8'hfe;
      17'd31973: data = 8'hfd;
      17'd31974: data = 8'hfc;
      17'd31975: data = 8'hfe;
      17'd31976: data = 8'hfd;
      17'd31977: data = 8'hf9;
      17'd31978: data = 8'hfd;
      17'd31979: data = 8'hfa;
      17'd31980: data = 8'hf9;
      17'd31981: data = 8'hfa;
      17'd31982: data = 8'hfc;
      17'd31983: data = 8'hfe;
      17'd31984: data = 8'h00;
      17'd31985: data = 8'h06;
      17'd31986: data = 8'h04;
      17'd31987: data = 8'h06;
      17'd31988: data = 8'h09;
      17'd31989: data = 8'h05;
      17'd31990: data = 8'h09;
      17'd31991: data = 8'h02;
      17'd31992: data = 8'h05;
      17'd31993: data = 8'h01;
      17'd31994: data = 8'h01;
      17'd31995: data = 8'h01;
      17'd31996: data = 8'hfc;
      17'd31997: data = 8'h02;
      17'd31998: data = 8'hfd;
      17'd31999: data = 8'hfa;
      17'd32000: data = 8'hfc;
      17'd32001: data = 8'hfe;
      17'd32002: data = 8'hfd;
      17'd32003: data = 8'hf5;
      17'd32004: data = 8'hfd;
      17'd32005: data = 8'h00;
      17'd32006: data = 8'hfd;
      17'd32007: data = 8'h00;
      17'd32008: data = 8'h01;
      17'd32009: data = 8'h04;
      17'd32010: data = 8'h01;
      17'd32011: data = 8'hfe;
      17'd32012: data = 8'h02;
      17'd32013: data = 8'hf4;
      17'd32014: data = 8'hf5;
      17'd32015: data = 8'hf6;
      17'd32016: data = 8'hed;
      17'd32017: data = 8'hed;
      17'd32018: data = 8'hf4;
      17'd32019: data = 8'hfc;
      17'd32020: data = 8'hf5;
      17'd32021: data = 8'hfa;
      17'd32022: data = 8'h02;
      17'd32023: data = 8'h06;
      17'd32024: data = 8'hf9;
      17'd32025: data = 8'hfc;
      17'd32026: data = 8'h00;
      17'd32027: data = 8'hf4;
      17'd32028: data = 8'hf5;
      17'd32029: data = 8'hef;
      17'd32030: data = 8'hfa;
      17'd32031: data = 8'hfd;
      17'd32032: data = 8'hec;
      17'd32033: data = 8'hf2;
      17'd32034: data = 8'hf6;
      17'd32035: data = 8'h04;
      17'd32036: data = 8'hfc;
      17'd32037: data = 8'he7;
      17'd32038: data = 8'hf4;
      17'd32039: data = 8'hf5;
      17'd32040: data = 8'hd2;
      17'd32041: data = 8'hc4;
      17'd32042: data = 8'hd8;
      17'd32043: data = 8'hd2;
      17'd32044: data = 8'hcb;
      17'd32045: data = 8'hd1;
      17'd32046: data = 8'hf4;
      17'd32047: data = 8'h11;
      17'd32048: data = 8'h05;
      17'd32049: data = 8'h29;
      17'd32050: data = 8'h4e;
      17'd32051: data = 8'h4f;
      17'd32052: data = 8'h52;
      17'd32053: data = 8'h4f;
      17'd32054: data = 8'h53;
      17'd32055: data = 8'h4a;
      17'd32056: data = 8'h3c;
      17'd32057: data = 8'h2d;
      17'd32058: data = 8'h1c;
      17'd32059: data = 8'h1b;
      17'd32060: data = 8'h0d;
      17'd32061: data = 8'hf6;
      17'd32062: data = 8'hec;
      17'd32063: data = 8'hf2;
      17'd32064: data = 8'hec;
      17'd32065: data = 8'hd1;
      17'd32066: data = 8'hd2;
      17'd32067: data = 8'he0;
      17'd32068: data = 8'hd6;
      17'd32069: data = 8'hc5;
      17'd32070: data = 8'hd3;
      17'd32071: data = 8'he4;
      17'd32072: data = 8'he4;
      17'd32073: data = 8'he4;
      17'd32074: data = 8'hed;
      17'd32075: data = 8'hfc;
      17'd32076: data = 8'hef;
      17'd32077: data = 8'hec;
      17'd32078: data = 8'heb;
      17'd32079: data = 8'he2;
      17'd32080: data = 8'he3;
      17'd32081: data = 8'hd5;
      17'd32082: data = 8'hcd;
      17'd32083: data = 8'hd1;
      17'd32084: data = 8'hd6;
      17'd32085: data = 8'hda;
      17'd32086: data = 8'hce;
      17'd32087: data = 8'hdc;
      17'd32088: data = 8'hef;
      17'd32089: data = 8'hed;
      17'd32090: data = 8'hef;
      17'd32091: data = 8'hfa;
      17'd32092: data = 8'h0d;
      17'd32093: data = 8'h12;
      17'd32094: data = 8'h13;
      17'd32095: data = 8'h22;
      17'd32096: data = 8'h2d;
      17'd32097: data = 8'h2f;
      17'd32098: data = 8'h29;
      17'd32099: data = 8'h2f;
      17'd32100: data = 8'h34;
      17'd32101: data = 8'h29;
      17'd32102: data = 8'h23;
      17'd32103: data = 8'h19;
      17'd32104: data = 8'h13;
      17'd32105: data = 8'h11;
      17'd32106: data = 8'h04;
      17'd32107: data = 8'h02;
      17'd32108: data = 8'h04;
      17'd32109: data = 8'h0a;
      17'd32110: data = 8'h11;
      17'd32111: data = 8'h0d;
      17'd32112: data = 8'h0e;
      17'd32113: data = 8'h1b;
      17'd32114: data = 8'h1c;
      17'd32115: data = 8'h15;
      17'd32116: data = 8'h1a;
      17'd32117: data = 8'h1e;
      17'd32118: data = 8'h1a;
      17'd32119: data = 8'h11;
      17'd32120: data = 8'h12;
      17'd32121: data = 8'h16;
      17'd32122: data = 8'h11;
      17'd32123: data = 8'h0c;
      17'd32124: data = 8'h09;
      17'd32125: data = 8'h0c;
      17'd32126: data = 8'h0a;
      17'd32127: data = 8'h01;
      17'd32128: data = 8'h00;
      17'd32129: data = 8'hfc;
      17'd32130: data = 8'h00;
      17'd32131: data = 8'hfc;
      17'd32132: data = 8'hf4;
      17'd32133: data = 8'hfd;
      17'd32134: data = 8'hfe;
      17'd32135: data = 8'hfd;
      17'd32136: data = 8'hfe;
      17'd32137: data = 8'h04;
      17'd32138: data = 8'h0e;
      17'd32139: data = 8'h0c;
      17'd32140: data = 8'h0a;
      17'd32141: data = 8'h12;
      17'd32142: data = 8'h13;
      17'd32143: data = 8'h0e;
      17'd32144: data = 8'h09;
      17'd32145: data = 8'h09;
      17'd32146: data = 8'h0a;
      17'd32147: data = 8'h06;
      17'd32148: data = 8'h01;
      17'd32149: data = 8'hfe;
      17'd32150: data = 8'h01;
      17'd32151: data = 8'h01;
      17'd32152: data = 8'hfa;
      17'd32153: data = 8'hfc;
      17'd32154: data = 8'h04;
      17'd32155: data = 8'h02;
      17'd32156: data = 8'hfe;
      17'd32157: data = 8'h05;
      17'd32158: data = 8'h0c;
      17'd32159: data = 8'h0a;
      17'd32160: data = 8'h02;
      17'd32161: data = 8'h02;
      17'd32162: data = 8'h05;
      17'd32163: data = 8'hf9;
      17'd32164: data = 8'hf6;
      17'd32165: data = 8'hf2;
      17'd32166: data = 8'hec;
      17'd32167: data = 8'he7;
      17'd32168: data = 8'he0;
      17'd32169: data = 8'he4;
      17'd32170: data = 8'he2;
      17'd32171: data = 8'he2;
      17'd32172: data = 8'he5;
      17'd32173: data = 8'he5;
      17'd32174: data = 8'he9;
      17'd32175: data = 8'hf1;
      17'd32176: data = 8'hed;
      17'd32177: data = 8'hec;
      17'd32178: data = 8'hf1;
      17'd32179: data = 8'hf1;
      17'd32180: data = 8'hec;
      17'd32181: data = 8'heb;
      17'd32182: data = 8'hed;
      17'd32183: data = 8'hed;
      17'd32184: data = 8'hec;
      17'd32185: data = 8'hed;
      17'd32186: data = 8'hf6;
      17'd32187: data = 8'hf2;
      17'd32188: data = 8'hf4;
      17'd32189: data = 8'hfa;
      17'd32190: data = 8'hf9;
      17'd32191: data = 8'hf9;
      17'd32192: data = 8'hf5;
      17'd32193: data = 8'hf9;
      17'd32194: data = 8'hf6;
      17'd32195: data = 8'hed;
      17'd32196: data = 8'hec;
      17'd32197: data = 8'hef;
      17'd32198: data = 8'hec;
      17'd32199: data = 8'hed;
      17'd32200: data = 8'hef;
      17'd32201: data = 8'hef;
      17'd32202: data = 8'hed;
      17'd32203: data = 8'heb;
      17'd32204: data = 8'he7;
      17'd32205: data = 8'hed;
      17'd32206: data = 8'hec;
      17'd32207: data = 8'he7;
      17'd32208: data = 8'hf1;
      17'd32209: data = 8'hf2;
      17'd32210: data = 8'hfa;
      17'd32211: data = 8'hfe;
      17'd32212: data = 8'h01;
      17'd32213: data = 8'h0a;
      17'd32214: data = 8'h04;
      17'd32215: data = 8'h0a;
      17'd32216: data = 8'h09;
      17'd32217: data = 8'h04;
      17'd32218: data = 8'h06;
      17'd32219: data = 8'h01;
      17'd32220: data = 8'hfe;
      17'd32221: data = 8'h00;
      17'd32222: data = 8'h06;
      17'd32223: data = 8'h02;
      17'd32224: data = 8'h01;
      17'd32225: data = 8'h02;
      17'd32226: data = 8'h05;
      17'd32227: data = 8'h02;
      17'd32228: data = 8'hfd;
      17'd32229: data = 8'h01;
      17'd32230: data = 8'hfa;
      17'd32231: data = 8'hf5;
      17'd32232: data = 8'hf1;
      17'd32233: data = 8'hef;
      17'd32234: data = 8'hed;
      17'd32235: data = 8'he5;
      17'd32236: data = 8'hed;
      17'd32237: data = 8'he9;
      17'd32238: data = 8'he9;
      17'd32239: data = 8'hfa;
      17'd32240: data = 8'hf5;
      17'd32241: data = 8'hf1;
      17'd32242: data = 8'hef;
      17'd32243: data = 8'he4;
      17'd32244: data = 8'hcd;
      17'd32245: data = 8'hbc;
      17'd32246: data = 8'hc5;
      17'd32247: data = 8'hc4;
      17'd32248: data = 8'hd1;
      17'd32249: data = 8'he4;
      17'd32250: data = 8'h04;
      17'd32251: data = 8'h27;
      17'd32252: data = 8'h3c;
      17'd32253: data = 8'h67;
      17'd32254: data = 8'h7d;
      17'd32255: data = 8'h7f;
      17'd32256: data = 8'h7f;
      17'd32257: data = 8'h7e;
      17'd32258: data = 8'h75;
      17'd32259: data = 8'h60;
      17'd32260: data = 8'h47;
      17'd32261: data = 8'h36;
      17'd32262: data = 8'h2d;
      17'd32263: data = 8'h19;
      17'd32264: data = 8'h09;
      17'd32265: data = 8'hfc;
      17'd32266: data = 8'hed;
      17'd32267: data = 8'he2;
      17'd32268: data = 8'hd2;
      17'd32269: data = 8'hcb;
      17'd32270: data = 8'hc6;
      17'd32271: data = 8'hbc;
      17'd32272: data = 8'hbc;
      17'd32273: data = 8'hbd;
      17'd32274: data = 8'hcd;
      17'd32275: data = 8'he3;
      17'd32276: data = 8'hed;
      17'd32277: data = 8'hfc;
      17'd32278: data = 8'h0a;
      17'd32279: data = 8'h0c;
      17'd32280: data = 8'h01;
      17'd32281: data = 8'hfd;
      17'd32282: data = 8'hfc;
      17'd32283: data = 8'hf2;
      17'd32284: data = 8'he2;
      17'd32285: data = 8'hda;
      17'd32286: data = 8'hdb;
      17'd32287: data = 8'hd5;
      17'd32288: data = 8'hd5;
      17'd32289: data = 8'hde;
      17'd32290: data = 8'heb;
      17'd32291: data = 8'hf9;
      17'd32292: data = 8'hfd;
      17'd32293: data = 8'h0a;
      17'd32294: data = 8'h1a;
      17'd32295: data = 8'h23;
      17'd32296: data = 8'h33;
      17'd32297: data = 8'h3a;
      17'd32298: data = 8'h46;
      17'd32299: data = 8'h52;
      17'd32300: data = 8'h52;
      17'd32301: data = 8'h4f;
      17'd32302: data = 8'h4b;
      17'd32303: data = 8'h43;
      17'd32304: data = 8'h33;
      17'd32305: data = 8'h1e;
      17'd32306: data = 8'h11;
      17'd32307: data = 8'h01;
      17'd32308: data = 8'hf1;
      17'd32309: data = 8'he7;
      17'd32310: data = 8'he7;
      17'd32311: data = 8'hed;
      17'd32312: data = 8'hf4;
      17'd32313: data = 8'hf5;
      17'd32314: data = 8'hfe;
      17'd32315: data = 8'h09;
      17'd32316: data = 8'h0a;
      17'd32317: data = 8'h0e;
      17'd32318: data = 8'h15;
      17'd32319: data = 8'h19;
      17'd32320: data = 8'h16;
      17'd32321: data = 8'h16;
      17'd32322: data = 8'h1b;
      17'd32323: data = 8'h1b;
      17'd32324: data = 8'h1e;
      17'd32325: data = 8'h1c;
      17'd32326: data = 8'h1a;
      17'd32327: data = 8'h15;
      17'd32328: data = 8'h0d;
      17'd32329: data = 8'h04;
      17'd32330: data = 8'hfc;
      17'd32331: data = 8'hf6;
      17'd32332: data = 8'hf9;
      17'd32333: data = 8'hfa;
      17'd32334: data = 8'hfc;
      17'd32335: data = 8'h01;
      17'd32336: data = 8'h0a;
      17'd32337: data = 8'h11;
      17'd32338: data = 8'h12;
      17'd32339: data = 8'h16;
      17'd32340: data = 8'h19;
      17'd32341: data = 8'h13;
      17'd32342: data = 8'h0d;
      17'd32343: data = 8'h09;
      17'd32344: data = 8'h01;
      17'd32345: data = 8'hfd;
      17'd32346: data = 8'hf6;
      17'd32347: data = 8'hf4;
      17'd32348: data = 8'hf2;
      17'd32349: data = 8'hed;
      17'd32350: data = 8'he5;
      17'd32351: data = 8'he5;
      17'd32352: data = 8'he7;
      17'd32353: data = 8'he3;
      17'd32354: data = 8'he2;
      17'd32355: data = 8'he3;
      17'd32356: data = 8'heb;
      17'd32357: data = 8'hef;
      17'd32358: data = 8'hf9;
      17'd32359: data = 8'h09;
      17'd32360: data = 8'h0a;
      17'd32361: data = 8'h09;
      17'd32362: data = 8'h13;
      17'd32363: data = 8'h05;
      17'd32364: data = 8'hf5;
      17'd32365: data = 8'h02;
      17'd32366: data = 8'hfc;
      17'd32367: data = 8'hed;
      17'd32368: data = 8'hf4;
      17'd32369: data = 8'hf9;
      17'd32370: data = 8'hf9;
      17'd32371: data = 8'hf1;
      17'd32372: data = 8'hf4;
      17'd32373: data = 8'h01;
      17'd32374: data = 8'hf6;
      17'd32375: data = 8'hf1;
      17'd32376: data = 8'hf6;
      17'd32377: data = 8'hed;
      17'd32378: data = 8'hed;
      17'd32379: data = 8'he9;
      17'd32380: data = 8'he7;
      17'd32381: data = 8'hec;
      17'd32382: data = 8'he9;
      17'd32383: data = 8'he7;
      17'd32384: data = 8'he4;
      17'd32385: data = 8'he7;
      17'd32386: data = 8'hed;
      17'd32387: data = 8'he2;
      17'd32388: data = 8'hde;
      17'd32389: data = 8'heb;
      17'd32390: data = 8'he4;
      17'd32391: data = 8'he4;
      17'd32392: data = 8'he7;
      17'd32393: data = 8'hf2;
      17'd32394: data = 8'hfc;
      17'd32395: data = 8'hf6;
      17'd32396: data = 8'hf9;
      17'd32397: data = 8'hfa;
      17'd32398: data = 8'hf4;
      17'd32399: data = 8'he9;
      17'd32400: data = 8'he5;
      17'd32401: data = 8'he4;
      17'd32402: data = 8'hde;
      17'd32403: data = 8'hd5;
      17'd32404: data = 8'hd6;
      17'd32405: data = 8'hd8;
      17'd32406: data = 8'hd6;
      17'd32407: data = 8'hd6;
      17'd32408: data = 8'hda;
      17'd32409: data = 8'he2;
      17'd32410: data = 8'he5;
      17'd32411: data = 8'he7;
      17'd32412: data = 8'hed;
      17'd32413: data = 8'hfa;
      17'd32414: data = 8'h00;
      17'd32415: data = 8'h05;
      17'd32416: data = 8'h0c;
      17'd32417: data = 8'h15;
      17'd32418: data = 8'h1c;
      17'd32419: data = 8'h1c;
      17'd32420: data = 8'h1b;
      17'd32421: data = 8'h1b;
      17'd32422: data = 8'h16;
      17'd32423: data = 8'h0e;
      17'd32424: data = 8'h06;
      17'd32425: data = 8'h02;
      17'd32426: data = 8'h01;
      17'd32427: data = 8'hfc;
      17'd32428: data = 8'hf9;
      17'd32429: data = 8'hfa;
      17'd32430: data = 8'hf6;
      17'd32431: data = 8'hf2;
      17'd32432: data = 8'hf2;
      17'd32433: data = 8'hec;
      17'd32434: data = 8'hf1;
      17'd32435: data = 8'hf2;
      17'd32436: data = 8'hef;
      17'd32437: data = 8'hfa;
      17'd32438: data = 8'hf9;
      17'd32439: data = 8'hfd;
      17'd32440: data = 8'h02;
      17'd32441: data = 8'h04;
      17'd32442: data = 8'h0a;
      17'd32443: data = 8'h04;
      17'd32444: data = 8'h06;
      17'd32445: data = 8'h0c;
      17'd32446: data = 8'h02;
      17'd32447: data = 8'h06;
      17'd32448: data = 8'h09;
      17'd32449: data = 8'h01;
      17'd32450: data = 8'h02;
      17'd32451: data = 8'hfd;
      17'd32452: data = 8'hfd;
      17'd32453: data = 8'h01;
      17'd32454: data = 8'hfc;
      17'd32455: data = 8'h01;
      17'd32456: data = 8'hf6;
      17'd32457: data = 8'hde;
      17'd32458: data = 8'hcb;
      17'd32459: data = 8'hb8;
      17'd32460: data = 8'hac;
      17'd32461: data = 8'hb1;
      17'd32462: data = 8'hc1;
      17'd32463: data = 8'hde;
      17'd32464: data = 8'h00;
      17'd32465: data = 8'h26;
      17'd32466: data = 8'h52;
      17'd32467: data = 8'h68;
      17'd32468: data = 8'h7f;
      17'd32469: data = 8'h7f;
      17'd32470: data = 8'h7f;
      17'd32471: data = 8'h7f;
      17'd32472: data = 8'h7f;
      17'd32473: data = 8'h6d;
      17'd32474: data = 8'h53;
      17'd32475: data = 8'h3a;
      17'd32476: data = 8'h26;
      17'd32477: data = 8'h12;
      17'd32478: data = 8'hfc;
      17'd32479: data = 8'he7;
      17'd32480: data = 8'hd3;
      17'd32481: data = 8'hc1;
      17'd32482: data = 8'hb9;
      17'd32483: data = 8'hb4;
      17'd32484: data = 8'hb5;
      17'd32485: data = 8'hbc;
      17'd32486: data = 8'hc9;
      17'd32487: data = 8'hd5;
      17'd32488: data = 8'he5;
      17'd32489: data = 8'hfd;
      17'd32490: data = 8'h19;
      17'd32491: data = 8'h29;
      17'd32492: data = 8'h33;
      17'd32493: data = 8'h2d;
      17'd32494: data = 8'h1f;
      17'd32495: data = 8'h0d;
      17'd32496: data = 8'hf6;
      17'd32497: data = 8'he9;
      17'd32498: data = 8'hdc;
      17'd32499: data = 8'hd2;
      17'd32500: data = 8'hc6;
      17'd32501: data = 8'hc4;
      17'd32502: data = 8'hc5;
      17'd32503: data = 8'hca;
      17'd32504: data = 8'hd3;
      17'd32505: data = 8'he0;
      17'd32506: data = 8'hf1;
      17'd32507: data = 8'hfe;
      17'd32508: data = 8'h0c;
      17'd32509: data = 8'h16;
      17'd32510: data = 8'h27;
      17'd32511: data = 8'h3a;
      17'd32512: data = 8'h47;
      17'd32513: data = 8'h4f;
      17'd32514: data = 8'h53;
      17'd32515: data = 8'h4d;
      17'd32516: data = 8'h3e;
      17'd32517: data = 8'h2c;
      17'd32518: data = 8'h16;
      17'd32519: data = 8'h02;
      17'd32520: data = 8'hef;
      17'd32521: data = 8'hdc;
      17'd32522: data = 8'hd1;
      17'd32523: data = 8'hca;
      17'd32524: data = 8'hca;
      17'd32525: data = 8'hd2;
      17'd32526: data = 8'he0;
      17'd32527: data = 8'hef;
      17'd32528: data = 8'hfd;
      17'd32529: data = 8'h06;
      17'd32530: data = 8'h12;
      17'd32531: data = 8'h1e;
      17'd32532: data = 8'h2c;
      17'd32533: data = 8'h34;
      17'd32534: data = 8'h39;
      17'd32535: data = 8'h3e;
      17'd32536: data = 8'h3d;
      17'd32537: data = 8'h39;
      17'd32538: data = 8'h31;
      17'd32539: data = 8'h27;
      17'd32540: data = 8'h1c;
      17'd32541: data = 8'h0e;
      17'd32542: data = 8'hfe;
      17'd32543: data = 8'hf2;
      17'd32544: data = 8'heb;
      17'd32545: data = 8'he3;
      17'd32546: data = 8'he3;
      17'd32547: data = 8'he5;
      17'd32548: data = 8'hf1;
      17'd32549: data = 8'hfd;
      17'd32550: data = 8'h02;
      17'd32551: data = 8'h09;
      17'd32552: data = 8'h0c;
      17'd32553: data = 8'h11;
      17'd32554: data = 8'h12;
      17'd32555: data = 8'h0c;
      17'd32556: data = 8'h06;
      17'd32557: data = 8'h04;
      17'd32558: data = 8'h00;
      17'd32559: data = 8'hfc;
      17'd32560: data = 8'hf9;
      17'd32561: data = 8'hf2;
      17'd32562: data = 8'he7;
      17'd32563: data = 8'he3;
      17'd32564: data = 8'he0;
      17'd32565: data = 8'hda;
      17'd32566: data = 8'hd8;
      17'd32567: data = 8'hda;
      17'd32568: data = 8'he0;
      17'd32569: data = 8'heb;
      17'd32570: data = 8'hf9;
      17'd32571: data = 8'h04;
      17'd32572: data = 8'h12;
      17'd32573: data = 8'h1c;
      17'd32574: data = 8'h26;
      17'd32575: data = 8'h29;
      17'd32576: data = 8'h26;
      17'd32577: data = 8'h22;
      17'd32578: data = 8'h1a;
      17'd32579: data = 8'h0d;
      17'd32580: data = 8'h01;
      17'd32581: data = 8'hf6;
      17'd32582: data = 8'hed;
      17'd32583: data = 8'he4;
      17'd32584: data = 8'hde;
      17'd32585: data = 8'hdc;
      17'd32586: data = 8'hd1;
      17'd32587: data = 8'hcb;
      17'd32588: data = 8'hd2;
      17'd32589: data = 8'hcb;
      17'd32590: data = 8'hcb;
      17'd32591: data = 8'hdb;
      17'd32592: data = 8'he2;
      17'd32593: data = 8'he4;
      17'd32594: data = 8'hf4;
      17'd32595: data = 8'h01;
      17'd32596: data = 8'h05;
      17'd32597: data = 8'h09;
      17'd32598: data = 8'h11;
      17'd32599: data = 8'h11;
      17'd32600: data = 8'h09;
      17'd32601: data = 8'h04;
      17'd32602: data = 8'h02;
      17'd32603: data = 8'hf9;
      17'd32604: data = 8'hf6;
      17'd32605: data = 8'hfd;
      17'd32606: data = 8'hf9;
      17'd32607: data = 8'hfc;
      17'd32608: data = 8'h00;
      17'd32609: data = 8'h01;
      17'd32610: data = 8'hfe;
      17'd32611: data = 8'hfe;
      17'd32612: data = 8'h00;
      17'd32613: data = 8'hf9;
      17'd32614: data = 8'hf1;
      17'd32615: data = 8'hec;
      17'd32616: data = 8'he5;
      17'd32617: data = 8'hde;
      17'd32618: data = 8'hd8;
      17'd32619: data = 8'hd6;
      17'd32620: data = 8'hd1;
      17'd32621: data = 8'hc9;
      17'd32622: data = 8'hc6;
      17'd32623: data = 8'hc9;
      17'd32624: data = 8'hce;
      17'd32625: data = 8'hd3;
      17'd32626: data = 8'he3;
      17'd32627: data = 8'hf2;
      17'd32628: data = 8'hfd;
      17'd32629: data = 8'h0d;
      17'd32630: data = 8'h1c;
      17'd32631: data = 8'h29;
      17'd32632: data = 8'h31;
      17'd32633: data = 8'h35;
      17'd32634: data = 8'h33;
      17'd32635: data = 8'h2b;
      17'd32636: data = 8'h24;
      17'd32637: data = 8'h16;
      17'd32638: data = 8'h0c;
      17'd32639: data = 8'h00;
      17'd32640: data = 8'hf5;
      17'd32641: data = 8'hef;
      17'd32642: data = 8'he5;
      17'd32643: data = 8'he2;
      17'd32644: data = 8'hdc;
      17'd32645: data = 8'hde;
      17'd32646: data = 8'he0;
      17'd32647: data = 8'he4;
      17'd32648: data = 8'he9;
      17'd32649: data = 8'hf1;
      17'd32650: data = 8'hf9;
      17'd32651: data = 8'hfc;
      17'd32652: data = 8'h06;
      17'd32653: data = 8'h0d;
      17'd32654: data = 8'h0e;
      17'd32655: data = 8'h12;
      17'd32656: data = 8'h13;
      17'd32657: data = 8'h11;
      17'd32658: data = 8'h09;
      17'd32659: data = 8'h02;
      17'd32660: data = 8'h01;
      17'd32661: data = 8'h00;
      17'd32662: data = 8'hf5;
      17'd32663: data = 8'hfa;
      17'd32664: data = 8'h01;
      17'd32665: data = 8'hfc;
      17'd32666: data = 8'h09;
      17'd32667: data = 8'h0d;
      17'd32668: data = 8'h13;
      17'd32669: data = 8'h1b;
      17'd32670: data = 8'h1c;
      17'd32671: data = 8'h2b;
      17'd32672: data = 8'h22;
      17'd32673: data = 8'h2c;
      17'd32674: data = 8'h31;
      17'd32675: data = 8'h2d;
      17'd32676: data = 8'h24;
      17'd32677: data = 8'h1a;
      17'd32678: data = 8'h02;
      17'd32679: data = 8'hc9;
      17'd32680: data = 8'hae;
      17'd32681: data = 8'h94;
      17'd32682: data = 8'h80;
      17'd32683: data = 8'h80;
      17'd32684: data = 8'h9f;
      17'd32685: data = 8'hb9;
      17'd32686: data = 8'hde;
      17'd32687: data = 8'h12;
      17'd32688: data = 8'h42;
      17'd32689: data = 8'h65;
      17'd32690: data = 8'h7f;
      17'd32691: data = 8'h7f;
      17'd32692: data = 8'h7f;
      17'd32693: data = 8'h7f;
      17'd32694: data = 8'h7f;
      17'd32695: data = 8'h7a;
      17'd32696: data = 8'h60;
      17'd32697: data = 8'h53;
      17'd32698: data = 8'h40;
      17'd32699: data = 8'h24;
      17'd32700: data = 8'h0c;
      17'd32701: data = 8'hed;
      17'd32702: data = 8'hd3;
      17'd32703: data = 8'hbc;
      17'd32704: data = 8'hae;
      17'd32705: data = 8'hb3;
      17'd32706: data = 8'hb9;
      17'd32707: data = 8'hc0;
      17'd32708: data = 8'hce;
      17'd32709: data = 8'he9;
      17'd32710: data = 8'hfe;
      17'd32711: data = 8'h0e;
      17'd32712: data = 8'h1f;
      17'd32713: data = 8'h24;
      17'd32714: data = 8'h19;
      17'd32715: data = 8'h06;
      17'd32716: data = 8'hf5;
      17'd32717: data = 8'hdc;
      17'd32718: data = 8'hc6;
      17'd32719: data = 8'hc1;
      17'd32720: data = 8'hbc;
      17'd32721: data = 8'hb9;
      17'd32722: data = 8'hbb;
      17'd32723: data = 8'hc0;
      17'd32724: data = 8'hc6;
      17'd32725: data = 8'hd3;
      17'd32726: data = 8'he2;
      17'd32727: data = 8'hf2;
      17'd32728: data = 8'h02;
      17'd32729: data = 8'h16;
      17'd32730: data = 8'h31;
      17'd32731: data = 8'h42;
      17'd32732: data = 8'h4e;
      17'd32733: data = 8'h56;
      17'd32734: data = 8'h5a;
      17'd32735: data = 8'h54;
      17'd32736: data = 8'h45;
      17'd32737: data = 8'h33;
      17'd32738: data = 8'h1b;
      17'd32739: data = 8'hfe;
      17'd32740: data = 8'heb;
      17'd32741: data = 8'hdb;
      17'd32742: data = 8'hcd;
      17'd32743: data = 8'hc6;
      17'd32744: data = 8'hc9;
      17'd32745: data = 8'hcd;
      17'd32746: data = 8'hd1;
      17'd32747: data = 8'hdb;
      17'd32748: data = 8'he4;
      17'd32749: data = 8'hef;
      17'd32750: data = 8'h01;
      17'd32751: data = 8'h12;
      17'd32752: data = 8'h1c;
      17'd32753: data = 8'h24;
      17'd32754: data = 8'h2c;
      17'd32755: data = 8'h33;
      17'd32756: data = 8'h31;
      17'd32757: data = 8'h2d;
      17'd32758: data = 8'h24;
      17'd32759: data = 8'h15;
      17'd32760: data = 8'h09;
      17'd32761: data = 8'hfc;
      17'd32762: data = 8'hed;
      17'd32763: data = 8'he5;
      17'd32764: data = 8'he5;
      17'd32765: data = 8'heb;
      17'd32766: data = 8'hf5;
      17'd32767: data = 8'h01;
      17'd32768: data = 8'h0a;
      17'd32769: data = 8'h12;
      17'd32770: data = 8'h1a;
      17'd32771: data = 8'h22;
      17'd32772: data = 8'h22;
      17'd32773: data = 8'h22;
      17'd32774: data = 8'h1e;
      17'd32775: data = 8'h1a;
      17'd32776: data = 8'h16;
      17'd32777: data = 8'h0e;
      17'd32778: data = 8'h04;
      17'd32779: data = 8'hfd;
      17'd32780: data = 8'hf2;
      17'd32781: data = 8'he7;
      17'd32782: data = 8'hdc;
      17'd32783: data = 8'hd5;
      17'd32784: data = 8'hd1;
      17'd32785: data = 8'hd2;
      17'd32786: data = 8'hdb;
      17'd32787: data = 8'he5;
      17'd32788: data = 8'hf4;
      17'd32789: data = 8'h04;
      17'd32790: data = 8'h15;
      17'd32791: data = 8'h1f;
      17'd32792: data = 8'h2b;
      17'd32793: data = 8'h2f;
      17'd32794: data = 8'h31;
      17'd32795: data = 8'h2b;
      17'd32796: data = 8'h26;
      17'd32797: data = 8'h1b;
      17'd32798: data = 8'h12;
      17'd32799: data = 8'h09;
      17'd32800: data = 8'hfd;
      17'd32801: data = 8'hf2;
      17'd32802: data = 8'he5;
      17'd32803: data = 8'hde;
      17'd32804: data = 8'hd5;
      17'd32805: data = 8'hd1;
      17'd32806: data = 8'hce;
      17'd32807: data = 8'hcd;
      17'd32808: data = 8'hd5;
      17'd32809: data = 8'hdc;
      17'd32810: data = 8'he5;
      17'd32811: data = 8'hef;
      17'd32812: data = 8'hf6;
      17'd32813: data = 8'h01;
      17'd32814: data = 8'h06;
      17'd32815: data = 8'h09;
      17'd32816: data = 8'h06;
      17'd32817: data = 8'hfd;
      17'd32818: data = 8'hf9;
      17'd32819: data = 8'hef;
      17'd32820: data = 8'he7;
      17'd32821: data = 8'heb;
      17'd32822: data = 8'he7;
      17'd32823: data = 8'he5;
      17'd32824: data = 8'heb;
      17'd32825: data = 8'hf4;
      17'd32826: data = 8'hfd;
      17'd32827: data = 8'h01;
      17'd32828: data = 8'h0d;
      17'd32829: data = 8'h16;
      17'd32830: data = 8'h1b;
      17'd32831: data = 8'h1f;
      17'd32832: data = 8'h22;
      17'd32833: data = 8'h22;
      17'd32834: data = 8'h19;
      17'd32835: data = 8'h12;
      17'd32836: data = 8'h02;
      17'd32837: data = 8'hf4;
      17'd32838: data = 8'he4;
      17'd32839: data = 8'hd6;
      17'd32840: data = 8'hce;
      17'd32841: data = 8'hc4;
      17'd32842: data = 8'hc0;
      17'd32843: data = 8'hc2;
      17'd32844: data = 8'hcd;
      17'd32845: data = 8'hd1;
      17'd32846: data = 8'hde;
      17'd32847: data = 8'hf1;
      17'd32848: data = 8'hfd;
      17'd32849: data = 8'h0a;
      17'd32850: data = 8'h19;
      17'd32851: data = 8'h1c;
      17'd32852: data = 8'h1e;
      17'd32853: data = 8'h24;
      17'd32854: data = 8'h23;
      17'd32855: data = 8'h22;
      17'd32856: data = 8'h1a;
      17'd32857: data = 8'h15;
      17'd32858: data = 8'h0a;
      17'd32859: data = 8'h01;
      17'd32860: data = 8'hfd;
      17'd32861: data = 8'hf4;
      17'd32862: data = 8'hec;
      17'd32863: data = 8'he9;
      17'd32864: data = 8'he4;
      17'd32865: data = 8'he2;
      17'd32866: data = 8'he3;
      17'd32867: data = 8'he5;
      17'd32868: data = 8'heb;
      17'd32869: data = 8'hec;
      17'd32870: data = 8'hef;
      17'd32871: data = 8'hf2;
      17'd32872: data = 8'hf2;
      17'd32873: data = 8'hfa;
      17'd32874: data = 8'hfa;
      17'd32875: data = 8'hfc;
      17'd32876: data = 8'h04;
      17'd32877: data = 8'hfd;
      17'd32878: data = 8'h09;
      17'd32879: data = 8'h09;
      17'd32880: data = 8'h09;
      17'd32881: data = 8'h01;
      17'd32882: data = 8'h06;
      17'd32883: data = 8'h0c;
      17'd32884: data = 8'hf5;
      17'd32885: data = 8'h13;
      17'd32886: data = 8'h00;
      17'd32887: data = 8'h06;
      17'd32888: data = 8'h13;
      17'd32889: data = 8'h09;
      17'd32890: data = 8'h19;
      17'd32891: data = 8'h0c;
      17'd32892: data = 8'h1b;
      17'd32893: data = 8'h1a;
      17'd32894: data = 8'h1b;
      17'd32895: data = 8'h26;
      17'd32896: data = 8'h24;
      17'd32897: data = 8'h1a;
      17'd32898: data = 8'h35;
      17'd32899: data = 8'h22;
      17'd32900: data = 8'h12;
      17'd32901: data = 8'h0e;
      17'd32902: data = 8'hd8;
      17'd32903: data = 8'hc2;
      17'd32904: data = 8'h95;
      17'd32905: data = 8'h8a;
      17'd32906: data = 8'h80;
      17'd32907: data = 8'h80;
      17'd32908: data = 8'ha4;
      17'd32909: data = 8'hc0;
      17'd32910: data = 8'hf6;
      17'd32911: data = 8'h2b;
      17'd32912: data = 8'h5f;
      17'd32913: data = 8'h7b;
      17'd32914: data = 8'h7f;
      17'd32915: data = 8'h7f;
      17'd32916: data = 8'h7f;
      17'd32917: data = 8'h7f;
      17'd32918: data = 8'h7f;
      17'd32919: data = 8'h64;
      17'd32920: data = 8'h4b;
      17'd32921: data = 8'h36;
      17'd32922: data = 8'h19;
      17'd32923: data = 8'h06;
      17'd32924: data = 8'he3;
      17'd32925: data = 8'hca;
      17'd32926: data = 8'hac;
      17'd32927: data = 8'ha4;
      17'd32928: data = 8'ha6;
      17'd32929: data = 8'hab;
      17'd32930: data = 8'hbc;
      17'd32931: data = 8'hd6;
      17'd32932: data = 8'hf1;
      17'd32933: data = 8'h0d;
      17'd32934: data = 8'h1c;
      17'd32935: data = 8'h22;
      17'd32936: data = 8'h22;
      17'd32937: data = 8'h13;
      17'd32938: data = 8'h04;
      17'd32939: data = 8'he5;
      17'd32940: data = 8'hd8;
      17'd32941: data = 8'hc9;
      17'd32942: data = 8'hbb;
      17'd32943: data = 8'hbb;
      17'd32944: data = 8'hb4;
      17'd32945: data = 8'hbd;
      17'd32946: data = 8'hc5;
      17'd32947: data = 8'hcd;
      17'd32948: data = 8'hde;
      17'd32949: data = 8'hec;
      17'd32950: data = 8'h02;
      17'd32951: data = 8'h13;
      17'd32952: data = 8'h27;
      17'd32953: data = 8'h42;
      17'd32954: data = 8'h4d;
      17'd32955: data = 8'h57;
      17'd32956: data = 8'h5b;
      17'd32957: data = 8'h53;
      17'd32958: data = 8'h42;
      17'd32959: data = 8'h26;
      17'd32960: data = 8'h0c;
      17'd32961: data = 8'hf2;
      17'd32962: data = 8'hda;
      17'd32963: data = 8'hc6;
      17'd32964: data = 8'hb4;
      17'd32965: data = 8'hb3;
      17'd32966: data = 8'hb9;
      17'd32967: data = 8'hc0;
      17'd32968: data = 8'hcd;
      17'd32969: data = 8'hda;
      17'd32970: data = 8'heb;
      17'd32971: data = 8'hfa;
      17'd32972: data = 8'h02;
      17'd32973: data = 8'h12;
      17'd32974: data = 8'h1e;
      17'd32975: data = 8'h29;
      17'd32976: data = 8'h31;
      17'd32977: data = 8'h34;
      17'd32978: data = 8'h33;
      17'd32979: data = 8'h27;
      17'd32980: data = 8'h1e;
      17'd32981: data = 8'h0e;
      17'd32982: data = 8'h00;
      17'd32983: data = 8'hf5;
      17'd32984: data = 8'hec;
      17'd32985: data = 8'he7;
      17'd32986: data = 8'heb;
      17'd32987: data = 8'hf2;
      17'd32988: data = 8'hfc;
      17'd32989: data = 8'h06;
      17'd32990: data = 8'h13;
      17'd32991: data = 8'h1e;
      17'd32992: data = 8'h23;
      17'd32993: data = 8'h24;
      17'd32994: data = 8'h24;
      17'd32995: data = 8'h1f;
      17'd32996: data = 8'h1b;
      17'd32997: data = 8'h12;
      17'd32998: data = 8'h0a;
      17'd32999: data = 8'h01;
      17'd33000: data = 8'hf4;
      17'd33001: data = 8'heb;
      17'd33002: data = 8'he0;
      17'd33003: data = 8'hd8;
      17'd33004: data = 8'hd2;
      17'd33005: data = 8'hd1;
      17'd33006: data = 8'hd5;
      17'd33007: data = 8'hde;
      17'd33008: data = 8'hed;
      17'd33009: data = 8'hfe;
      17'd33010: data = 8'h0e;
      17'd33011: data = 8'h1c;
      17'd33012: data = 8'h2c;
      17'd33013: data = 8'h33;
      17'd33014: data = 8'h35;
      17'd33015: data = 8'h33;
      17'd33016: data = 8'h2b;
      17'd33017: data = 8'h1f;
      17'd33018: data = 8'h13;
      17'd33019: data = 8'h09;
      17'd33020: data = 8'h00;
      17'd33021: data = 8'hf5;
      17'd33022: data = 8'he7;
      17'd33023: data = 8'he2;
      17'd33024: data = 8'hdb;
      17'd33025: data = 8'hd6;
      17'd33026: data = 8'hd6;
      17'd33027: data = 8'hd6;
      17'd33028: data = 8'hdc;
      17'd33029: data = 8'he5;
      17'd33030: data = 8'hef;
      17'd33031: data = 8'hfd;
      17'd33032: data = 8'h04;
      17'd33033: data = 8'h0c;
      17'd33034: data = 8'h0e;
      17'd33035: data = 8'h11;
      17'd33036: data = 8'h0e;
      17'd33037: data = 8'h06;
      17'd33038: data = 8'h01;
      17'd33039: data = 8'hf9;
      17'd33040: data = 8'hf4;
      17'd33041: data = 8'hf1;
      17'd33042: data = 8'hec;
      17'd33043: data = 8'hf1;
      17'd33044: data = 8'hf4;
      17'd33045: data = 8'hf5;
      17'd33046: data = 8'hfa;
      17'd33047: data = 8'h00;
      17'd33048: data = 8'h05;
      17'd33049: data = 8'h09;
      17'd33050: data = 8'h0e;
      17'd33051: data = 8'h12;
      17'd33052: data = 8'h13;
      17'd33053: data = 8'h12;
      17'd33054: data = 8'h05;
      17'd33055: data = 8'h02;
      17'd33056: data = 8'hf5;
      17'd33057: data = 8'he0;
      17'd33058: data = 8'hd3;
      17'd33059: data = 8'hd1;
      17'd33060: data = 8'hc2;
      17'd33061: data = 8'hbd;
      17'd33062: data = 8'hc6;
      17'd33063: data = 8'hca;
      17'd33064: data = 8'hd1;
      17'd33065: data = 8'he4;
      17'd33066: data = 8'hf9;
      17'd33067: data = 8'hf2;
      17'd33068: data = 8'h06;
      17'd33069: data = 8'h16;
      17'd33070: data = 8'h19;
      17'd33071: data = 8'h23;
      17'd33072: data = 8'h2c;
      17'd33073: data = 8'h2f;
      17'd33074: data = 8'h27;
      17'd33075: data = 8'h2f;
      17'd33076: data = 8'h27;
      17'd33077: data = 8'h1c;
      17'd33078: data = 8'h12;
      17'd33079: data = 8'h0d;
      17'd33080: data = 8'hfd;
      17'd33081: data = 8'hf1;
      17'd33082: data = 8'hec;
      17'd33083: data = 8'he3;
      17'd33084: data = 8'he3;
      17'd33085: data = 8'he0;
      17'd33086: data = 8'he7;
      17'd33087: data = 8'he4;
      17'd33088: data = 8'he9;
      17'd33089: data = 8'heb;
      17'd33090: data = 8'hed;
      17'd33091: data = 8'hec;
      17'd33092: data = 8'hf1;
      17'd33093: data = 8'hf6;
      17'd33094: data = 8'hfc;
      17'd33095: data = 8'hfe;
      17'd33096: data = 8'h04;
      17'd33097: data = 8'h0a;
      17'd33098: data = 8'h09;
      17'd33099: data = 8'h0e;
      17'd33100: data = 8'h11;
      17'd33101: data = 8'h0a;
      17'd33102: data = 8'h05;
      17'd33103: data = 8'h09;
      17'd33104: data = 8'h00;
      17'd33105: data = 8'hfa;
      17'd33106: data = 8'hf5;
      17'd33107: data = 8'hed;
      17'd33108: data = 8'hec;
      17'd33109: data = 8'he7;
      17'd33110: data = 8'he9;
      17'd33111: data = 8'he7;
      17'd33112: data = 8'hec;
      17'd33113: data = 8'hec;
      17'd33114: data = 8'hf6;
      17'd33115: data = 8'h04;
      17'd33116: data = 8'h0a;
      17'd33117: data = 8'h15;
      17'd33118: data = 8'h1c;
      17'd33119: data = 8'h23;
      17'd33120: data = 8'h1e;
      17'd33121: data = 8'h1f;
      17'd33122: data = 8'h22;
      17'd33123: data = 8'h12;
      17'd33124: data = 8'h0e;
      17'd33125: data = 8'h0e;
      17'd33126: data = 8'h00;
      17'd33127: data = 8'hfe;
      17'd33128: data = 8'hfd;
      17'd33129: data = 8'hfe;
      17'd33130: data = 8'hfa;
      17'd33131: data = 8'hf1;
      17'd33132: data = 8'hf6;
      17'd33133: data = 8'hf6;
      17'd33134: data = 8'he2;
      17'd33135: data = 8'he2;
      17'd33136: data = 8'hde;
      17'd33137: data = 8'hb9;
      17'd33138: data = 8'hae;
      17'd33139: data = 8'hac;
      17'd33140: data = 8'haa;
      17'd33141: data = 8'ha4;
      17'd33142: data = 8'hcd;
      17'd33143: data = 8'hfa;
      17'd33144: data = 8'h0a;
      17'd33145: data = 8'h39;
      17'd33146: data = 8'h65;
      17'd33147: data = 8'h72;
      17'd33148: data = 8'h7f;
      17'd33149: data = 8'h7f;
      17'd33150: data = 8'h7f;
      17'd33151: data = 8'h7f;
      17'd33152: data = 8'h7b;
      17'd33153: data = 8'h68;
      17'd33154: data = 8'h45;
      17'd33155: data = 8'h2c;
      17'd33156: data = 8'h16;
      17'd33157: data = 8'hf5;
      17'd33158: data = 8'hda;
      17'd33159: data = 8'hc0;
      17'd33160: data = 8'ha6;
      17'd33161: data = 8'h94;
      17'd33162: data = 8'h97;
      17'd33163: data = 8'h9d;
      17'd33164: data = 8'haa;
      17'd33165: data = 8'hb9;
      17'd33166: data = 8'hcd;
      17'd33167: data = 8'he2;
      17'd33168: data = 8'hef;
      17'd33169: data = 8'hfa;
      17'd33170: data = 8'hfe;
      17'd33171: data = 8'hfc;
      17'd33172: data = 8'hfa;
      17'd33173: data = 8'hf2;
      17'd33174: data = 8'hed;
      17'd33175: data = 8'heb;
      17'd33176: data = 8'he7;
      17'd33177: data = 8'heb;
      17'd33178: data = 8'hec;
      17'd33179: data = 8'hf1;
      17'd33180: data = 8'hf9;
      17'd33181: data = 8'hfd;
      17'd33182: data = 8'h06;
      17'd33183: data = 8'h11;
      17'd33184: data = 8'h19;
      17'd33185: data = 8'h24;
      17'd33186: data = 8'h2d;
      17'd33187: data = 8'h36;
      17'd33188: data = 8'h3a;
      17'd33189: data = 8'h36;
      17'd33190: data = 8'h31;
      17'd33191: data = 8'h1f;
      17'd33192: data = 8'h0e;
      17'd33193: data = 8'hf9;
      17'd33194: data = 8'hde;
      17'd33195: data = 8'hcb;
      17'd33196: data = 8'hbd;
      17'd33197: data = 8'hb5;
      17'd33198: data = 8'hb0;
      17'd33199: data = 8'hb0;
      17'd33200: data = 8'hb8;
      17'd33201: data = 8'hc2;
      17'd33202: data = 8'hd2;
      17'd33203: data = 8'he2;
      17'd33204: data = 8'hf5;
      17'd33205: data = 8'h05;
      17'd33206: data = 8'h16;
      17'd33207: data = 8'h29;
      17'd33208: data = 8'h39;
      17'd33209: data = 8'h40;
      17'd33210: data = 8'h46;
      17'd33211: data = 8'h4b;
      17'd33212: data = 8'h45;
      17'd33213: data = 8'h3d;
      17'd33214: data = 8'h35;
      17'd33215: data = 8'h27;
      17'd33216: data = 8'h19;
      17'd33217: data = 8'h0d;
      17'd33218: data = 8'h04;
      17'd33219: data = 8'hfd;
      17'd33220: data = 8'hfe;
      17'd33221: data = 8'h00;
      17'd33222: data = 8'hfe;
      17'd33223: data = 8'hfd;
      17'd33224: data = 8'h00;
      17'd33225: data = 8'h01;
      17'd33226: data = 8'h00;
      17'd33227: data = 8'hfe;
      17'd33228: data = 8'hf9;
      17'd33229: data = 8'hf4;
      17'd33230: data = 8'hf1;
      17'd33231: data = 8'hed;
      17'd33232: data = 8'he9;
      17'd33233: data = 8'he5;
      17'd33234: data = 8'he3;
      17'd33235: data = 8'he0;
      17'd33236: data = 8'he0;
      17'd33237: data = 8'he2;
      17'd33238: data = 8'he7;
      17'd33239: data = 8'hf1;
      17'd33240: data = 8'hfa;
      17'd33241: data = 8'h09;
      17'd33242: data = 8'h19;
      17'd33243: data = 8'h26;
      17'd33244: data = 8'h33;
      17'd33245: data = 8'h3a;
      17'd33246: data = 8'h3e;
      17'd33247: data = 8'h3e;
      17'd33248: data = 8'h3d;
      17'd33249: data = 8'h3a;
      17'd33250: data = 8'h2f;
      17'd33251: data = 8'h23;
      17'd33252: data = 8'h15;
      17'd33253: data = 8'h09;
      17'd33254: data = 8'hfc;
      17'd33255: data = 8'hf1;
      17'd33256: data = 8'he5;
      17'd33257: data = 8'hdb;
      17'd33258: data = 8'hd3;
      17'd33259: data = 8'hcd;
      17'd33260: data = 8'hcd;
      17'd33261: data = 8'hd2;
      17'd33262: data = 8'hd6;
      17'd33263: data = 8'hdb;
      17'd33264: data = 8'he4;
      17'd33265: data = 8'hed;
      17'd33266: data = 8'hf4;
      17'd33267: data = 8'hf6;
      17'd33268: data = 8'hfa;
      17'd33269: data = 8'hfa;
      17'd33270: data = 8'hf9;
      17'd33271: data = 8'hf5;
      17'd33272: data = 8'hf6;
      17'd33273: data = 8'hf5;
      17'd33274: data = 8'hf4;
      17'd33275: data = 8'hf5;
      17'd33276: data = 8'hfa;
      17'd33277: data = 8'h01;
      17'd33278: data = 8'h09;
      17'd33279: data = 8'h0d;
      17'd33280: data = 8'h15;
      17'd33281: data = 8'h1a;
      17'd33282: data = 8'h1e;
      17'd33283: data = 8'h22;
      17'd33284: data = 8'h23;
      17'd33285: data = 8'h23;
      17'd33286: data = 8'h1e;
      17'd33287: data = 8'h16;
      17'd33288: data = 8'h11;
      17'd33289: data = 8'h06;
      17'd33290: data = 8'hf5;
      17'd33291: data = 8'he3;
      17'd33292: data = 8'hca;
      17'd33293: data = 8'hb4;
      17'd33294: data = 8'hae;
      17'd33295: data = 8'hab;
      17'd33296: data = 8'ha6;
      17'd33297: data = 8'hb0;
      17'd33298: data = 8'hc1;
      17'd33299: data = 8'hcb;
      17'd33300: data = 8'he0;
      17'd33301: data = 8'hfa;
      17'd33302: data = 8'h0a;
      17'd33303: data = 8'h15;
      17'd33304: data = 8'h2d;
      17'd33305: data = 8'h39;
      17'd33306: data = 8'h3c;
      17'd33307: data = 8'h46;
      17'd33308: data = 8'h4a;
      17'd33309: data = 8'h40;
      17'd33310: data = 8'h3e;
      17'd33311: data = 8'h3a;
      17'd33312: data = 8'h26;
      17'd33313: data = 8'h13;
      17'd33314: data = 8'h06;
      17'd33315: data = 8'hf9;
      17'd33316: data = 8'he9;
      17'd33317: data = 8'he9;
      17'd33318: data = 8'he3;
      17'd33319: data = 8'hdb;
      17'd33320: data = 8'hde;
      17'd33321: data = 8'hde;
      17'd33322: data = 8'hde;
      17'd33323: data = 8'he4;
      17'd33324: data = 8'he2;
      17'd33325: data = 8'he3;
      17'd33326: data = 8'he4;
      17'd33327: data = 8'heb;
      17'd33328: data = 8'hf4;
      17'd33329: data = 8'hf9;
      17'd33330: data = 8'hfd;
      17'd33331: data = 8'hfe;
      17'd33332: data = 8'h02;
      17'd33333: data = 8'h09;
      17'd33334: data = 8'h06;
      17'd33335: data = 8'h0c;
      17'd33336: data = 8'h0e;
      17'd33337: data = 8'h04;
      17'd33338: data = 8'h11;
      17'd33339: data = 8'h11;
      17'd33340: data = 8'h0c;
      17'd33341: data = 8'h09;
      17'd33342: data = 8'h05;
      17'd33343: data = 8'h01;
      17'd33344: data = 8'hf6;
      17'd33345: data = 8'hf5;
      17'd33346: data = 8'hec;
      17'd33347: data = 8'hec;
      17'd33348: data = 8'hf1;
      17'd33349: data = 8'hf2;
      17'd33350: data = 8'hf4;
      17'd33351: data = 8'h06;
      17'd33352: data = 8'h06;
      17'd33353: data = 8'h06;
      17'd33354: data = 8'h0e;
      17'd33355: data = 8'h16;
      17'd33356: data = 8'h0d;
      17'd33357: data = 8'h12;
      17'd33358: data = 8'h16;
      17'd33359: data = 8'h01;
      17'd33360: data = 8'hfc;
      17'd33361: data = 8'h0d;
      17'd33362: data = 8'hf6;
      17'd33363: data = 8'heb;
      17'd33364: data = 8'h00;
      17'd33365: data = 8'hde;
      17'd33366: data = 8'hfe;
      17'd33367: data = 8'hed;
      17'd33368: data = 8'hfd;
      17'd33369: data = 8'h00;
      17'd33370: data = 8'hec;
      17'd33371: data = 8'h01;
      17'd33372: data = 8'he3;
      17'd33373: data = 8'heb;
      17'd33374: data = 8'hda;
      17'd33375: data = 8'hbd;
      17'd33376: data = 8'hcb;
      17'd33377: data = 8'hbc;
      17'd33378: data = 8'hc6;
      17'd33379: data = 8'hf6;
      17'd33380: data = 8'h02;
      17'd33381: data = 8'h2d;
      17'd33382: data = 8'h40;
      17'd33383: data = 8'h53;
      17'd33384: data = 8'h60;
      17'd33385: data = 8'h63;
      17'd33386: data = 8'h77;
      17'd33387: data = 8'h67;
      17'd33388: data = 8'h63;
      17'd33389: data = 8'h68;
      17'd33390: data = 8'h4a;
      17'd33391: data = 8'h3a;
      17'd33392: data = 8'h2b;
      17'd33393: data = 8'h0d;
      17'd33394: data = 8'hfc;
      17'd33395: data = 8'he3;
      17'd33396: data = 8'hd8;
      17'd33397: data = 8'hc0;
      17'd33398: data = 8'hb4;
      17'd33399: data = 8'hbc;
      17'd33400: data = 8'hbd;
      17'd33401: data = 8'hce;
      17'd33402: data = 8'hdb;
      17'd33403: data = 8'he7;
      17'd33404: data = 8'hf4;
      17'd33405: data = 8'hf5;
      17'd33406: data = 8'hf2;
      17'd33407: data = 8'hf6;
      17'd33408: data = 8'heb;
      17'd33409: data = 8'heb;
      17'd33410: data = 8'heb;
      17'd33411: data = 8'he4;
      17'd33412: data = 8'he5;
      17'd33413: data = 8'he5;
      17'd33414: data = 8'heb;
      17'd33415: data = 8'he5;
      17'd33416: data = 8'heb;
      17'd33417: data = 8'hf5;
      17'd33418: data = 8'hfd;
      17'd33419: data = 8'h06;
      17'd33420: data = 8'h12;
      17'd33421: data = 8'h1a;
      17'd33422: data = 8'h23;
      17'd33423: data = 8'h2b;
      17'd33424: data = 8'h34;
      17'd33425: data = 8'h35;
      17'd33426: data = 8'h31;
      17'd33427: data = 8'h23;
      17'd33428: data = 8'h13;
      17'd33429: data = 8'h05;
      17'd33430: data = 8'hf4;
      17'd33431: data = 8'heb;
      17'd33432: data = 8'hde;
      17'd33433: data = 8'hd8;
      17'd33434: data = 8'hd8;
      17'd33435: data = 8'hd2;
      17'd33436: data = 8'hd6;
      17'd33437: data = 8'hd6;
      17'd33438: data = 8'hdb;
      17'd33439: data = 8'he4;
      17'd33440: data = 8'hec;
      17'd33441: data = 8'hfc;
      17'd33442: data = 8'h02;
      17'd33443: data = 8'h0e;
      17'd33444: data = 8'h19;
      17'd33445: data = 8'h1c;
      17'd33446: data = 8'h27;
      17'd33447: data = 8'h2b;
      17'd33448: data = 8'h29;
      17'd33449: data = 8'h26;
      17'd33450: data = 8'h1e;
      17'd33451: data = 8'h1a;
      17'd33452: data = 8'h11;
      17'd33453: data = 8'h0d;
      17'd33454: data = 8'h0c;
      17'd33455: data = 8'h0a;
      17'd33456: data = 8'h0e;
      17'd33457: data = 8'h13;
      17'd33458: data = 8'h19;
      17'd33459: data = 8'h19;
      17'd33460: data = 8'h1a;
      17'd33461: data = 8'h1b;
      17'd33462: data = 8'h1b;
      17'd33463: data = 8'h1c;
      17'd33464: data = 8'h1a;
      17'd33465: data = 8'h13;
      17'd33466: data = 8'h0c;
      17'd33467: data = 8'h01;
      17'd33468: data = 8'hf4;
      17'd33469: data = 8'he9;
      17'd33470: data = 8'hdc;
      17'd33471: data = 8'hd6;
      17'd33472: data = 8'hcd;
      17'd33473: data = 8'hca;
      17'd33474: data = 8'hcb;
      17'd33475: data = 8'hd1;
      17'd33476: data = 8'hdc;
      17'd33477: data = 8'he9;
      17'd33478: data = 8'hf6;
      17'd33479: data = 8'h06;
      17'd33480: data = 8'h15;
      17'd33481: data = 8'h1b;
      17'd33482: data = 8'h24;
      17'd33483: data = 8'h2c;
      17'd33484: data = 8'h2d;
      17'd33485: data = 8'h2d;
      17'd33486: data = 8'h2d;
      17'd33487: data = 8'h29;
      17'd33488: data = 8'h1f;
      17'd33489: data = 8'h19;
      17'd33490: data = 8'h0e;
      17'd33491: data = 8'h05;
      17'd33492: data = 8'hfd;
      17'd33493: data = 8'hf5;
      17'd33494: data = 8'hed;
      17'd33495: data = 8'he7;
      17'd33496: data = 8'he5;
      17'd33497: data = 8'he5;
      17'd33498: data = 8'he7;
      17'd33499: data = 8'heb;
      17'd33500: data = 8'heb;
      17'd33501: data = 8'hec;
      17'd33502: data = 8'hec;
      17'd33503: data = 8'he9;
      17'd33504: data = 8'he7;
      17'd33505: data = 8'he4;
      17'd33506: data = 8'he3;
      17'd33507: data = 8'he3;
      17'd33508: data = 8'he4;
      17'd33509: data = 8'he5;
      17'd33510: data = 8'he7;
      17'd33511: data = 8'heb;
      17'd33512: data = 8'hf1;
      17'd33513: data = 8'hf6;
      17'd33514: data = 8'hfe;
      17'd33515: data = 8'h05;
      17'd33516: data = 8'h0e;
      17'd33517: data = 8'h1a;
      17'd33518: data = 8'h22;
      17'd33519: data = 8'h23;
      17'd33520: data = 8'h23;
      17'd33521: data = 8'h22;
      17'd33522: data = 8'h1a;
      17'd33523: data = 8'h13;
      17'd33524: data = 8'h0c;
      17'd33525: data = 8'h00;
      17'd33526: data = 8'hf4;
      17'd33527: data = 8'heb;
      17'd33528: data = 8'he4;
      17'd33529: data = 8'hda;
      17'd33530: data = 8'hda;
      17'd33531: data = 8'hdb;
      17'd33532: data = 8'hd8;
      17'd33533: data = 8'hdb;
      17'd33534: data = 8'he4;
      17'd33535: data = 8'heb;
      17'd33536: data = 8'hec;
      17'd33537: data = 8'hf4;
      17'd33538: data = 8'hfd;
      17'd33539: data = 8'hfc;
      17'd33540: data = 8'h00;
      17'd33541: data = 8'h09;
      17'd33542: data = 8'h05;
      17'd33543: data = 8'h05;
      17'd33544: data = 8'h0a;
      17'd33545: data = 8'h0a;
      17'd33546: data = 8'h06;
      17'd33547: data = 8'h06;
      17'd33548: data = 8'h06;
      17'd33549: data = 8'h06;
      17'd33550: data = 8'h09;
      17'd33551: data = 8'h09;
      17'd33552: data = 8'h05;
      17'd33553: data = 8'h01;
      17'd33554: data = 8'h00;
      17'd33555: data = 8'hfd;
      17'd33556: data = 8'hfd;
      17'd33557: data = 8'hfa;
      17'd33558: data = 8'hf5;
      17'd33559: data = 8'hf5;
      17'd33560: data = 8'hed;
      17'd33561: data = 8'hef;
      17'd33562: data = 8'hf1;
      17'd33563: data = 8'hed;
      17'd33564: data = 8'heb;
      17'd33565: data = 8'hef;
      17'd33566: data = 8'hef;
      17'd33567: data = 8'hf2;
      17'd33568: data = 8'hfa;
      17'd33569: data = 8'hfd;
      17'd33570: data = 8'hfe;
      17'd33571: data = 8'h00;
      17'd33572: data = 8'h06;
      17'd33573: data = 8'h05;
      17'd33574: data = 8'h02;
      17'd33575: data = 8'h01;
      17'd33576: data = 8'hfa;
      17'd33577: data = 8'hef;
      17'd33578: data = 8'hf6;
      17'd33579: data = 8'hed;
      17'd33580: data = 8'he9;
      17'd33581: data = 8'hef;
      17'd33582: data = 8'hef;
      17'd33583: data = 8'hfc;
      17'd33584: data = 8'hfd;
      17'd33585: data = 8'h0c;
      17'd33586: data = 8'h13;
      17'd33587: data = 8'h11;
      17'd33588: data = 8'h15;
      17'd33589: data = 8'h1c;
      17'd33590: data = 8'h15;
      17'd33591: data = 8'h0e;
      17'd33592: data = 8'h0a;
      17'd33593: data = 8'h0c;
      17'd33594: data = 8'h01;
      17'd33595: data = 8'hf9;
      17'd33596: data = 8'h01;
      17'd33597: data = 8'hf4;
      17'd33598: data = 8'hf6;
      17'd33599: data = 8'h01;
      17'd33600: data = 8'h01;
      17'd33601: data = 8'h02;
      17'd33602: data = 8'h06;
      17'd33603: data = 8'hfe;
      17'd33604: data = 8'hfa;
      17'd33605: data = 8'he9;
      17'd33606: data = 8'he7;
      17'd33607: data = 8'he2;
      17'd33608: data = 8'hc2;
      17'd33609: data = 8'hbc;
      17'd33610: data = 8'ha6;
      17'd33611: data = 8'hb4;
      17'd33612: data = 8'hb0;
      17'd33613: data = 8'hc5;
      17'd33614: data = 8'hf5;
      17'd33615: data = 8'h05;
      17'd33616: data = 8'h2d;
      17'd33617: data = 8'h4e;
      17'd33618: data = 8'h5f;
      17'd33619: data = 8'h6c;
      17'd33620: data = 8'h74;
      17'd33621: data = 8'h7e;
      17'd33622: data = 8'h77;
      17'd33623: data = 8'h72;
      17'd33624: data = 8'h74;
      17'd33625: data = 8'h4b;
      17'd33626: data = 8'h3c;
      17'd33627: data = 8'h27;
      17'd33628: data = 8'h06;
      17'd33629: data = 8'hf1;
      17'd33630: data = 8'hde;
      17'd33631: data = 8'hd2;
      17'd33632: data = 8'hb9;
      17'd33633: data = 8'hb5;
      17'd33634: data = 8'hc2;
      17'd33635: data = 8'hc5;
      17'd33636: data = 8'hd6;
      17'd33637: data = 8'he4;
      17'd33638: data = 8'hf1;
      17'd33639: data = 8'hf9;
      17'd33640: data = 8'hfd;
      17'd33641: data = 8'hfd;
      17'd33642: data = 8'hf4;
      17'd33643: data = 8'hf2;
      17'd33644: data = 8'hed;
      17'd33645: data = 8'heb;
      17'd33646: data = 8'he7;
      17'd33647: data = 8'he4;
      17'd33648: data = 8'hdc;
      17'd33649: data = 8'hda;
      17'd33650: data = 8'hdb;
      17'd33651: data = 8'he5;
      17'd33652: data = 8'hef;
      17'd33653: data = 8'hf6;
      17'd33654: data = 8'h06;
      17'd33655: data = 8'h13;
      17'd33656: data = 8'h1e;
      17'd33657: data = 8'h2b;
      17'd33658: data = 8'h35;
      17'd33659: data = 8'h36;
      17'd33660: data = 8'h35;
      17'd33661: data = 8'h2f;
      17'd33662: data = 8'h22;
      17'd33663: data = 8'h0d;
      17'd33664: data = 8'hfe;
      17'd33665: data = 8'hec;
      17'd33666: data = 8'hde;
      17'd33667: data = 8'hd8;
      17'd33668: data = 8'hd5;
      17'd33669: data = 8'hd1;
      17'd33670: data = 8'hca;
      17'd33671: data = 8'hcd;
      17'd33672: data = 8'hd2;
      17'd33673: data = 8'hdc;
      17'd33674: data = 8'heb;
      17'd33675: data = 8'hf6;
      17'd33676: data = 8'h04;
      17'd33677: data = 8'h0a;
      17'd33678: data = 8'h15;
      17'd33679: data = 8'h1e;
      17'd33680: data = 8'h1f;
      17'd33681: data = 8'h22;
      17'd33682: data = 8'h1e;
      17'd33683: data = 8'h1a;
      17'd33684: data = 8'h12;
      17'd33685: data = 8'h0d;
      17'd33686: data = 8'h09;
      17'd33687: data = 8'h04;
      17'd33688: data = 8'h06;
      17'd33689: data = 8'h0c;
      17'd33690: data = 8'h12;
      17'd33691: data = 8'h19;
      17'd33692: data = 8'h1c;
      17'd33693: data = 8'h1e;
      17'd33694: data = 8'h22;
      17'd33695: data = 8'h26;
      17'd33696: data = 8'h27;
      17'd33697: data = 8'h23;
      17'd33698: data = 8'h1c;
      17'd33699: data = 8'h16;
      17'd33700: data = 8'h0a;
      17'd33701: data = 8'h00;
      17'd33702: data = 8'hf5;
      17'd33703: data = 8'he3;
      17'd33704: data = 8'hd5;
      17'd33705: data = 8'hcb;
      17'd33706: data = 8'hc6;
      17'd33707: data = 8'hc9;
      17'd33708: data = 8'hcb;
      17'd33709: data = 8'hd3;
      17'd33710: data = 8'hdc;
      17'd33711: data = 8'hed;
      17'd33712: data = 8'hfd;
      17'd33713: data = 8'h06;
      17'd33714: data = 8'h11;
      17'd33715: data = 8'h1b;
      17'd33716: data = 8'h1f;
      17'd33717: data = 8'h26;
      17'd33718: data = 8'h27;
      17'd33719: data = 8'h27;
      17'd33720: data = 8'h26;
      17'd33721: data = 8'h22;
      17'd33722: data = 8'h1e;
      17'd33723: data = 8'h16;
      17'd33724: data = 8'h11;
      17'd33725: data = 8'h06;
      17'd33726: data = 8'h00;
      17'd33727: data = 8'hfd;
      17'd33728: data = 8'hfc;
      17'd33729: data = 8'hfc;
      17'd33730: data = 8'hf9;
      17'd33731: data = 8'hf9;
      17'd33732: data = 8'hf6;
      17'd33733: data = 8'hf5;
      17'd33734: data = 8'hf9;
      17'd33735: data = 8'hf4;
      17'd33736: data = 8'hed;
      17'd33737: data = 8'he7;
      17'd33738: data = 8'he4;
      17'd33739: data = 8'hde;
      17'd33740: data = 8'hdc;
      17'd33741: data = 8'hdc;
      17'd33742: data = 8'hda;
      17'd33743: data = 8'hda;
      17'd33744: data = 8'hde;
      17'd33745: data = 8'he7;
      17'd33746: data = 8'hed;
      17'd33747: data = 8'hf5;
      17'd33748: data = 8'hf6;
      17'd33749: data = 8'hfc;
      17'd33750: data = 8'h0a;
      17'd33751: data = 8'h13;
      17'd33752: data = 8'h1b;
      17'd33753: data = 8'h24;
      17'd33754: data = 8'h26;
      17'd33755: data = 8'h27;
      17'd33756: data = 8'h27;
      17'd33757: data = 8'h1f;
      17'd33758: data = 8'h19;
      17'd33759: data = 8'h0c;
      17'd33760: data = 8'h01;
      17'd33761: data = 8'hfc;
      17'd33762: data = 8'hf9;
      17'd33763: data = 8'hf4;
      17'd33764: data = 8'he5;
      17'd33765: data = 8'he3;
      17'd33766: data = 8'he3;
      17'd33767: data = 8'he2;
      17'd33768: data = 8'he0;
      17'd33769: data = 8'hde;
      17'd33770: data = 8'hda;
      17'd33771: data = 8'hdb;
      17'd33772: data = 8'he2;
      17'd33773: data = 8'he7;
      17'd33774: data = 8'hec;
      17'd33775: data = 8'hef;
      17'd33776: data = 8'hf2;
      17'd33777: data = 8'hf9;
      17'd33778: data = 8'h04;
      17'd33779: data = 8'h0a;
      17'd33780: data = 8'h0a;
      17'd33781: data = 8'h0a;
      17'd33782: data = 8'h13;
      17'd33783: data = 8'h1a;
      17'd33784: data = 8'h1e;
      17'd33785: data = 8'h23;
      17'd33786: data = 8'h1e;
      17'd33787: data = 8'h19;
      17'd33788: data = 8'h13;
      17'd33789: data = 8'h0d;
      17'd33790: data = 8'h04;
      17'd33791: data = 8'h01;
      17'd33792: data = 8'hf2;
      17'd33793: data = 8'he7;
      17'd33794: data = 8'he7;
      17'd33795: data = 8'he4;
      17'd33796: data = 8'he3;
      17'd33797: data = 8'hdc;
      17'd33798: data = 8'hde;
      17'd33799: data = 8'he0;
      17'd33800: data = 8'he4;
      17'd33801: data = 8'hef;
      17'd33802: data = 8'hf2;
      17'd33803: data = 8'hf4;
      17'd33804: data = 8'hfd;
      17'd33805: data = 8'hfc;
      17'd33806: data = 8'h01;
      17'd33807: data = 8'h0c;
      17'd33808: data = 8'h04;
      17'd33809: data = 8'h04;
      17'd33810: data = 8'h01;
      17'd33811: data = 8'h01;
      17'd33812: data = 8'h06;
      17'd33813: data = 8'hfc;
      17'd33814: data = 8'h06;
      17'd33815: data = 8'h06;
      17'd33816: data = 8'h04;
      17'd33817: data = 8'h0c;
      17'd33818: data = 8'h0d;
      17'd33819: data = 8'h19;
      17'd33820: data = 8'hfe;
      17'd33821: data = 8'h12;
      17'd33822: data = 8'h1c;
      17'd33823: data = 8'h01;
      17'd33824: data = 8'h24;
      17'd33825: data = 8'h12;
      17'd33826: data = 8'h05;
      17'd33827: data = 8'h16;
      17'd33828: data = 8'h0d;
      17'd33829: data = 8'h19;
      17'd33830: data = 8'h09;
      17'd33831: data = 8'h05;
      17'd33832: data = 8'h01;
      17'd33833: data = 8'he0;
      17'd33834: data = 8'hf2;
      17'd33835: data = 8'he2;
      17'd33836: data = 8'hc2;
      17'd33837: data = 8'hcd;
      17'd33838: data = 8'hab;
      17'd33839: data = 8'h9b;
      17'd33840: data = 8'h97;
      17'd33841: data = 8'h9b;
      17'd33842: data = 8'hb0;
      17'd33843: data = 8'hc1;
      17'd33844: data = 8'hfd;
      17'd33845: data = 8'h16;
      17'd33846: data = 8'h31;
      17'd33847: data = 8'h5f;
      17'd33848: data = 8'h64;
      17'd33849: data = 8'h72;
      17'd33850: data = 8'h7f;
      17'd33851: data = 8'h7f;
      17'd33852: data = 8'h7f;
      17'd33853: data = 8'h7f;
      17'd33854: data = 8'h7b;
      17'd33855: data = 8'h5b;
      17'd33856: data = 8'h3d;
      17'd33857: data = 8'h34;
      17'd33858: data = 8'h0d;
      17'd33859: data = 8'hf2;
      17'd33860: data = 8'he2;
      17'd33861: data = 8'hc9;
      17'd33862: data = 8'hbd;
      17'd33863: data = 8'hc0;
      17'd33864: data = 8'hd1;
      17'd33865: data = 8'hd1;
      17'd33866: data = 8'hde;
      17'd33867: data = 8'heb;
      17'd33868: data = 8'he9;
      17'd33869: data = 8'heb;
      17'd33870: data = 8'heb;
      17'd33871: data = 8'he5;
      17'd33872: data = 8'he0;
      17'd33873: data = 8'hde;
      17'd33874: data = 8'hdc;
      17'd33875: data = 8'hd1;
      17'd33876: data = 8'hc9;
      17'd33877: data = 8'hc5;
      17'd33878: data = 8'hc0;
      17'd33879: data = 8'hca;
      17'd33880: data = 8'hd3;
      17'd33881: data = 8'he0;
      17'd33882: data = 8'hf1;
      17'd33883: data = 8'hfc;
      17'd33884: data = 8'h12;
      17'd33885: data = 8'h24;
      17'd33886: data = 8'h36;
      17'd33887: data = 8'h47;
      17'd33888: data = 8'h4f;
      17'd33889: data = 8'h54;
      17'd33890: data = 8'h4b;
      17'd33891: data = 8'h3e;
      17'd33892: data = 8'h2d;
      17'd33893: data = 8'h16;
      17'd33894: data = 8'h05;
      17'd33895: data = 8'hf6;
      17'd33896: data = 8'he7;
      17'd33897: data = 8'hdb;
      17'd33898: data = 8'hce;
      17'd33899: data = 8'hca;
      17'd33900: data = 8'hc4;
      17'd33901: data = 8'hca;
      17'd33902: data = 8'hd5;
      17'd33903: data = 8'hde;
      17'd33904: data = 8'hed;
      17'd33905: data = 8'hf9;
      17'd33906: data = 8'h05;
      17'd33907: data = 8'h0e;
      17'd33908: data = 8'h15;
      17'd33909: data = 8'h1a;
      17'd33910: data = 8'h16;
      17'd33911: data = 8'h12;
      17'd33912: data = 8'h0e;
      17'd33913: data = 8'h05;
      17'd33914: data = 8'hfe;
      17'd33915: data = 8'hfc;
      17'd33916: data = 8'hfa;
      17'd33917: data = 8'h00;
      17'd33918: data = 8'h05;
      17'd33919: data = 8'h0c;
      17'd33920: data = 8'h12;
      17'd33921: data = 8'h16;
      17'd33922: data = 8'h22;
      17'd33923: data = 8'h2b;
      17'd33924: data = 8'h34;
      17'd33925: data = 8'h3a;
      17'd33926: data = 8'h3c;
      17'd33927: data = 8'h3a;
      17'd33928: data = 8'h34;
      17'd33929: data = 8'h2c;
      17'd33930: data = 8'h22;
      17'd33931: data = 8'h11;
      17'd33932: data = 8'h04;
      17'd33933: data = 8'hf5;
      17'd33934: data = 8'he7;
      17'd33935: data = 8'hdc;
      17'd33936: data = 8'hd1;
      17'd33937: data = 8'hcd;
      17'd33938: data = 8'hcd;
      17'd33939: data = 8'hd1;
      17'd33940: data = 8'hd6;
      17'd33941: data = 8'hdc;
      17'd33942: data = 8'he5;
      17'd33943: data = 8'hef;
      17'd33944: data = 8'hf9;
      17'd33945: data = 8'h06;
      17'd33946: data = 8'h0e;
      17'd33947: data = 8'h16;
      17'd33948: data = 8'h1a;
      17'd33949: data = 8'h16;
      17'd33950: data = 8'h15;
      17'd33951: data = 8'h0e;
      17'd33952: data = 8'h0d;
      17'd33953: data = 8'h09;
      17'd33954: data = 8'h04;
      17'd33955: data = 8'h04;
      17'd33956: data = 8'h01;
      17'd33957: data = 8'h04;
      17'd33958: data = 8'h05;
      17'd33959: data = 8'h09;
      17'd33960: data = 8'h0e;
      17'd33961: data = 8'h13;
      17'd33962: data = 8'h15;
      17'd33963: data = 8'h15;
      17'd33964: data = 8'h12;
      17'd33965: data = 8'h0d;
      17'd33966: data = 8'h09;
      17'd33967: data = 8'h04;
      17'd33968: data = 8'hfc;
      17'd33969: data = 8'hef;
      17'd33970: data = 8'he4;
      17'd33971: data = 8'hdb;
      17'd33972: data = 8'hd6;
      17'd33973: data = 8'hc9;
      17'd33974: data = 8'hbc;
      17'd33975: data = 8'hbb;
      17'd33976: data = 8'hbb;
      17'd33977: data = 8'hc0;
      17'd33978: data = 8'hce;
      17'd33979: data = 8'he0;
      17'd33980: data = 8'heb;
      17'd33981: data = 8'hfa;
      17'd33982: data = 8'h0a;
      17'd33983: data = 8'h15;
      17'd33984: data = 8'h1b;
      17'd33985: data = 8'h1f;
      17'd33986: data = 8'h22;
      17'd33987: data = 8'h1f;
      17'd33988: data = 8'h24;
      17'd33989: data = 8'h23;
      17'd33990: data = 8'h16;
      17'd33991: data = 8'h13;
      17'd33992: data = 8'h0e;
      17'd33993: data = 8'h04;
      17'd33994: data = 8'hf9;
      17'd33995: data = 8'hf1;
      17'd33996: data = 8'he9;
      17'd33997: data = 8'hde;
      17'd33998: data = 8'he3;
      17'd33999: data = 8'he7;
      17'd34000: data = 8'he2;
      17'd34001: data = 8'hde;
      17'd34002: data = 8'hde;
      17'd34003: data = 8'he0;
      17'd34004: data = 8'he0;
      17'd34005: data = 8'he7;
      17'd34006: data = 8'he9;
      17'd34007: data = 8'he7;
      17'd34008: data = 8'hf1;
      17'd34009: data = 8'hf9;
      17'd34010: data = 8'hfe;
      17'd34011: data = 8'h05;
      17'd34012: data = 8'h0d;
      17'd34013: data = 8'h13;
      17'd34014: data = 8'h19;
      17'd34015: data = 8'h22;
      17'd34016: data = 8'h24;
      17'd34017: data = 8'h1f;
      17'd34018: data = 8'h1a;
      17'd34019: data = 8'h16;
      17'd34020: data = 8'h12;
      17'd34021: data = 8'h09;
      17'd34022: data = 8'h00;
      17'd34023: data = 8'hf4;
      17'd34024: data = 8'heb;
      17'd34025: data = 8'he3;
      17'd34026: data = 8'he2;
      17'd34027: data = 8'hdc;
      17'd34028: data = 8'hd8;
      17'd34029: data = 8'hd6;
      17'd34030: data = 8'hdb;
      17'd34031: data = 8'he4;
      17'd34032: data = 8'heb;
      17'd34033: data = 8'hf5;
      17'd34034: data = 8'hf4;
      17'd34035: data = 8'h00;
      17'd34036: data = 8'h05;
      17'd34037: data = 8'h04;
      17'd34038: data = 8'h0a;
      17'd34039: data = 8'h05;
      17'd34040: data = 8'h06;
      17'd34041: data = 8'hfe;
      17'd34042: data = 8'h01;
      17'd34043: data = 8'h09;
      17'd34044: data = 8'hfc;
      17'd34045: data = 8'h01;
      17'd34046: data = 8'h0d;
      17'd34047: data = 8'h00;
      17'd34048: data = 8'h15;
      17'd34049: data = 8'h12;
      17'd34050: data = 8'h1b;
      17'd34051: data = 8'h1c;
      17'd34052: data = 8'h06;
      17'd34053: data = 8'h2f;
      17'd34054: data = 8'h0a;
      17'd34055: data = 8'h1b;
      17'd34056: data = 8'h3c;
      17'd34057: data = 8'h1b;
      17'd34058: data = 8'h0e;
      17'd34059: data = 8'hf2;
      17'd34060: data = 8'hdc;
      17'd34061: data = 8'hc1;
      17'd34062: data = 8'h99;
      17'd34063: data = 8'hca;
      17'd34064: data = 8'he0;
      17'd34065: data = 8'hd1;
      17'd34066: data = 8'h04;
      17'd34067: data = 8'hf6;
      17'd34068: data = 8'hef;
      17'd34069: data = 8'hf1;
      17'd34070: data = 8'hf5;
      17'd34071: data = 8'h05;
      17'd34072: data = 8'h02;
      17'd34073: data = 8'h27;
      17'd34074: data = 8'h31;
      17'd34075: data = 8'h22;
      17'd34076: data = 8'h46;
      17'd34077: data = 8'h43;
      17'd34078: data = 8'h2d;
      17'd34079: data = 8'h34;
      17'd34080: data = 8'h2d;
      17'd34081: data = 8'h2f;
      17'd34082: data = 8'h16;
      17'd34083: data = 8'h2b;
      17'd34084: data = 8'h39;
      17'd34085: data = 8'h27;
      17'd34086: data = 8'h39;
      17'd34087: data = 8'h24;
      17'd34088: data = 8'h13;
      17'd34089: data = 8'h09;
      17'd34090: data = 8'hfe;
      17'd34091: data = 8'h04;
      17'd34092: data = 8'h01;
      17'd34093: data = 8'hfe;
      17'd34094: data = 8'hf1;
      17'd34095: data = 8'hd8;
      17'd34096: data = 8'hd6;
      17'd34097: data = 8'hc9;
      17'd34098: data = 8'hbd;
      17'd34099: data = 8'hc4;
      17'd34100: data = 8'hc4;
      17'd34101: data = 8'hcd;
      17'd34102: data = 8'hd1;
      17'd34103: data = 8'hd8;
      17'd34104: data = 8'hda;
      17'd34105: data = 8'hda;
      17'd34106: data = 8'hda;
      17'd34107: data = 8'hde;
      17'd34108: data = 8'he9;
      17'd34109: data = 8'hf5;
      17'd34110: data = 8'hfc;
      17'd34111: data = 8'h05;
      17'd34112: data = 8'h19;
      17'd34113: data = 8'h22;
      17'd34114: data = 8'h23;
      17'd34115: data = 8'h22;
      17'd34116: data = 8'h1a;
      17'd34117: data = 8'h13;
      17'd34118: data = 8'h13;
      17'd34119: data = 8'h16;
      17'd34120: data = 8'h1a;
      17'd34121: data = 8'h19;
      17'd34122: data = 8'h16;
      17'd34123: data = 8'h13;
      17'd34124: data = 8'h0d;
      17'd34125: data = 8'h0e;
      17'd34126: data = 8'h00;
      17'd34127: data = 8'hf6;
      17'd34128: data = 8'hf6;
      17'd34129: data = 8'hf5;
      17'd34130: data = 8'hf4;
      17'd34131: data = 8'hf2;
      17'd34132: data = 8'hf9;
      17'd34133: data = 8'hf4;
      17'd34134: data = 8'hf1;
      17'd34135: data = 8'hf4;
      17'd34136: data = 8'hf1;
      17'd34137: data = 8'hed;
      17'd34138: data = 8'hed;
      17'd34139: data = 8'hf2;
      17'd34140: data = 8'hfc;
      17'd34141: data = 8'h05;
      17'd34142: data = 8'h0a;
      17'd34143: data = 8'h0d;
      17'd34144: data = 8'h0d;
      17'd34145: data = 8'h13;
      17'd34146: data = 8'h13;
      17'd34147: data = 8'h15;
      17'd34148: data = 8'h1a;
      17'd34149: data = 8'h1a;
      17'd34150: data = 8'h1e;
      17'd34151: data = 8'h22;
      17'd34152: data = 8'h22;
      17'd34153: data = 8'h1b;
      17'd34154: data = 8'h11;
      17'd34155: data = 8'h0a;
      17'd34156: data = 8'h05;
      17'd34157: data = 8'h04;
      17'd34158: data = 8'h09;
      17'd34159: data = 8'h02;
      17'd34160: data = 8'h02;
      17'd34161: data = 8'h06;
      17'd34162: data = 8'h06;
      17'd34163: data = 8'h05;
      17'd34164: data = 8'h01;
      17'd34165: data = 8'h02;
      17'd34166: data = 8'hfe;
      17'd34167: data = 8'hfe;
      17'd34168: data = 8'h04;
      17'd34169: data = 8'h04;
      17'd34170: data = 8'h02;
      17'd34171: data = 8'h02;
      17'd34172: data = 8'h00;
      17'd34173: data = 8'hfd;
      17'd34174: data = 8'hf5;
      17'd34175: data = 8'hf1;
      17'd34176: data = 8'hed;
      17'd34177: data = 8'hf1;
      17'd34178: data = 8'hfa;
      17'd34179: data = 8'hfc;
      17'd34180: data = 8'hfe;
      17'd34181: data = 8'h01;
      17'd34182: data = 8'h04;
      17'd34183: data = 8'h02;
      17'd34184: data = 8'h02;
      17'd34185: data = 8'h06;
      17'd34186: data = 8'h04;
      17'd34187: data = 8'h01;
      17'd34188: data = 8'h04;
      17'd34189: data = 8'h05;
      17'd34190: data = 8'h05;
      17'd34191: data = 8'h02;
      17'd34192: data = 8'hfd;
      17'd34193: data = 8'hfa;
      17'd34194: data = 8'hf5;
      17'd34195: data = 8'hf4;
      17'd34196: data = 8'hfc;
      17'd34197: data = 8'hf5;
      17'd34198: data = 8'hed;
      17'd34199: data = 8'he9;
      17'd34200: data = 8'hf1;
      17'd34201: data = 8'hf2;
      17'd34202: data = 8'heb;
      17'd34203: data = 8'hed;
      17'd34204: data = 8'hef;
      17'd34205: data = 8'heb;
      17'd34206: data = 8'hf5;
      17'd34207: data = 8'hfd;
      17'd34208: data = 8'hf4;
      17'd34209: data = 8'hef;
      17'd34210: data = 8'hf4;
      17'd34211: data = 8'hfc;
      17'd34212: data = 8'hfc;
      17'd34213: data = 8'hfa;
      17'd34214: data = 8'hf6;
      17'd34215: data = 8'hf2;
      17'd34216: data = 8'hf9;
      17'd34217: data = 8'h04;
      17'd34218: data = 8'hfe;
      17'd34219: data = 8'hfa;
      17'd34220: data = 8'hfd;
      17'd34221: data = 8'hfc;
      17'd34222: data = 8'hfa;
      17'd34223: data = 8'hfc;
      17'd34224: data = 8'hf9;
      17'd34225: data = 8'hf1;
      17'd34226: data = 8'hf4;
      17'd34227: data = 8'hfd;
      17'd34228: data = 8'hfa;
      17'd34229: data = 8'hed;
      17'd34230: data = 8'he9;
      17'd34231: data = 8'he5;
      17'd34232: data = 8'he7;
      17'd34233: data = 8'hed;
      17'd34234: data = 8'hec;
      17'd34235: data = 8'hf1;
      17'd34236: data = 8'hfc;
      17'd34237: data = 8'hfa;
      17'd34238: data = 8'h01;
      17'd34239: data = 8'h04;
      17'd34240: data = 8'h01;
      17'd34241: data = 8'h09;
      17'd34242: data = 8'h02;
      17'd34243: data = 8'h02;
      17'd34244: data = 8'h0d;
      17'd34245: data = 8'h09;
      17'd34246: data = 8'h01;
      17'd34247: data = 8'h05;
      17'd34248: data = 8'hfe;
      17'd34249: data = 8'hf9;
      17'd34250: data = 8'hfe;
      17'd34251: data = 8'hf4;
      17'd34252: data = 8'hef;
      17'd34253: data = 8'hf1;
      17'd34254: data = 8'hf1;
      17'd34255: data = 8'hf6;
      17'd34256: data = 8'hf9;
      17'd34257: data = 8'hf2;
      17'd34258: data = 8'hef;
      17'd34259: data = 8'hec;
      17'd34260: data = 8'hf9;
      17'd34261: data = 8'hfc;
      17'd34262: data = 8'hf1;
      17'd34263: data = 8'hf2;
      17'd34264: data = 8'hfa;
      17'd34265: data = 8'h00;
      17'd34266: data = 8'h00;
      17'd34267: data = 8'h09;
      17'd34268: data = 8'h0a;
      17'd34269: data = 8'h00;
      17'd34270: data = 8'h0c;
      17'd34271: data = 8'h06;
      17'd34272: data = 8'h04;
      17'd34273: data = 8'h0c;
      17'd34274: data = 8'h04;
      17'd34275: data = 8'h06;
      17'd34276: data = 8'h06;
      17'd34277: data = 8'h0e;
      17'd34278: data = 8'h0e;
      17'd34279: data = 8'hfe;
      17'd34280: data = 8'h0a;
      17'd34281: data = 8'h19;
      17'd34282: data = 8'h00;
      17'd34283: data = 8'h0e;
      17'd34284: data = 8'h0d;
      17'd34285: data = 8'h0a;
      17'd34286: data = 8'h11;
      17'd34287: data = 8'h02;
      17'd34288: data = 8'h12;
      17'd34289: data = 8'hf6;
      17'd34290: data = 8'h00;
      17'd34291: data = 8'h06;
      17'd34292: data = 8'he9;
      17'd34293: data = 8'hfa;
      17'd34294: data = 8'hf4;
      17'd34295: data = 8'he7;
      17'd34296: data = 8'he3;
      17'd34297: data = 8'hc2;
      17'd34298: data = 8'hc4;
      17'd34299: data = 8'hc2;
      17'd34300: data = 8'hdb;
      17'd34301: data = 8'hf2;
      17'd34302: data = 8'hf2;
      17'd34303: data = 8'h16;
      17'd34304: data = 8'h24;
      17'd34305: data = 8'h2d;
      17'd34306: data = 8'h3d;
      17'd34307: data = 8'h45;
      17'd34308: data = 8'h36;
      17'd34309: data = 8'h29;
      17'd34310: data = 8'h42;
      17'd34311: data = 8'h3e;
      17'd34312: data = 8'h27;
      17'd34313: data = 8'h23;
      17'd34314: data = 8'h1f;
      17'd34315: data = 8'h13;
      17'd34316: data = 8'h01;
      17'd34317: data = 8'hfe;
      17'd34318: data = 8'hed;
      17'd34319: data = 8'he3;
      17'd34320: data = 8'hf6;
      17'd34321: data = 8'hfc;
      17'd34322: data = 8'h00;
      17'd34323: data = 8'h05;
      17'd34324: data = 8'h02;
      17'd34325: data = 8'hf9;
      17'd34326: data = 8'hed;
      17'd34327: data = 8'hf9;
      17'd34328: data = 8'hf1;
      17'd34329: data = 8'he5;
      17'd34330: data = 8'hed;
      17'd34331: data = 8'hed;
      17'd34332: data = 8'heb;
      17'd34333: data = 8'hed;
      17'd34334: data = 8'hf1;
      17'd34335: data = 8'hdc;
      17'd34336: data = 8'hd1;
      17'd34337: data = 8'hd8;
      17'd34338: data = 8'hdb;
      17'd34339: data = 8'he2;
      17'd34340: data = 8'hec;
      17'd34341: data = 8'hf2;
      17'd34342: data = 8'hf6;
      17'd34343: data = 8'h01;
      17'd34344: data = 8'h0e;
      17'd34345: data = 8'h09;
      17'd34346: data = 8'h04;
      17'd34347: data = 8'h05;
      17'd34348: data = 8'h09;
      17'd34349: data = 8'h0e;
      17'd34350: data = 8'h13;
      17'd34351: data = 8'h15;
      17'd34352: data = 8'h0c;
      17'd34353: data = 8'h0c;
      17'd34354: data = 8'h0c;
      17'd34355: data = 8'h02;
      17'd34356: data = 8'hfe;
      17'd34357: data = 8'hfa;
      17'd34358: data = 8'hfa;
      17'd34359: data = 8'hfd;
      17'd34360: data = 8'h05;
      17'd34361: data = 8'h0e;
      17'd34362: data = 8'h06;
      17'd34363: data = 8'h09;
      17'd34364: data = 8'h06;
      17'd34365: data = 8'h06;
      17'd34366: data = 8'h0c;
      17'd34367: data = 8'h06;
      17'd34368: data = 8'h05;
      17'd34369: data = 8'h06;
      17'd34370: data = 8'h0c;
      17'd34371: data = 8'h0d;
      17'd34372: data = 8'h0c;
      17'd34373: data = 8'h09;
      17'd34374: data = 8'h00;
      17'd34375: data = 8'h00;
      17'd34376: data = 8'h02;
      17'd34377: data = 8'h02;
      17'd34378: data = 8'h05;
      17'd34379: data = 8'h04;
      17'd34380: data = 8'h05;
      17'd34381: data = 8'h09;
      17'd34382: data = 8'h09;
      17'd34383: data = 8'h0a;
      17'd34384: data = 8'h01;
      17'd34385: data = 8'h00;
      17'd34386: data = 8'h02;
      17'd34387: data = 8'h01;
      17'd34388: data = 8'h06;
      17'd34389: data = 8'h09;
      17'd34390: data = 8'h06;
      17'd34391: data = 8'h04;
      17'd34392: data = 8'h06;
      17'd34393: data = 8'h0a;
      17'd34394: data = 8'h04;
      17'd34395: data = 8'h02;
      17'd34396: data = 8'h02;
      17'd34397: data = 8'h05;
      17'd34398: data = 8'h0c;
      17'd34399: data = 8'h0e;
      17'd34400: data = 8'h11;
      17'd34401: data = 8'h0c;
      17'd34402: data = 8'h09;
      17'd34403: data = 8'h0d;
      17'd34404: data = 8'h06;
      17'd34405: data = 8'h04;
      17'd34406: data = 8'h02;
      17'd34407: data = 8'hfd;
      17'd34408: data = 8'h00;
      17'd34409: data = 8'h01;
      17'd34410: data = 8'hfe;
      17'd34411: data = 8'hfa;
      17'd34412: data = 8'hf4;
      17'd34413: data = 8'hf4;
      17'd34414: data = 8'hf2;
      17'd34415: data = 8'hf4;
      17'd34416: data = 8'hf5;
      17'd34417: data = 8'hf4;
      17'd34418: data = 8'hf5;
      17'd34419: data = 8'hf6;
      17'd34420: data = 8'hf6;
      17'd34421: data = 8'hf5;
      17'd34422: data = 8'hf4;
      17'd34423: data = 8'hf1;
      17'd34424: data = 8'hf4;
      17'd34425: data = 8'hf6;
      17'd34426: data = 8'hf1;
      17'd34427: data = 8'hef;
      17'd34428: data = 8'hf5;
      17'd34429: data = 8'hf6;
      17'd34430: data = 8'hfa;
      17'd34431: data = 8'hfa;
      17'd34432: data = 8'hfd;
      17'd34433: data = 8'hfc;
      17'd34434: data = 8'hfc;
      17'd34435: data = 8'h04;
      17'd34436: data = 8'h05;
      17'd34437: data = 8'hfe;
      17'd34438: data = 8'h00;
      17'd34439: data = 8'h04;
      17'd34440: data = 8'h00;
      17'd34441: data = 8'hfd;
      17'd34442: data = 8'hfc;
      17'd34443: data = 8'hfa;
      17'd34444: data = 8'hf6;
      17'd34445: data = 8'hfa;
      17'd34446: data = 8'hfa;
      17'd34447: data = 8'hf9;
      17'd34448: data = 8'hf6;
      17'd34449: data = 8'hf5;
      17'd34450: data = 8'hf4;
      17'd34451: data = 8'hf2;
      17'd34452: data = 8'hf1;
      17'd34453: data = 8'hef;
      17'd34454: data = 8'heb;
      17'd34455: data = 8'heb;
      17'd34456: data = 8'hed;
      17'd34457: data = 8'heb;
      17'd34458: data = 8'he9;
      17'd34459: data = 8'he7;
      17'd34460: data = 8'he9;
      17'd34461: data = 8'he9;
      17'd34462: data = 8'heb;
      17'd34463: data = 8'hef;
      17'd34464: data = 8'hed;
      17'd34465: data = 8'hef;
      17'd34466: data = 8'hf5;
      17'd34467: data = 8'hf9;
      17'd34468: data = 8'hfe;
      17'd34469: data = 8'hfe;
      17'd34470: data = 8'h00;
      17'd34471: data = 8'h02;
      17'd34472: data = 8'h05;
      17'd34473: data = 8'h06;
      17'd34474: data = 8'h05;
      17'd34475: data = 8'h02;
      17'd34476: data = 8'h00;
      17'd34477: data = 8'hfc;
      17'd34478: data = 8'hfc;
      17'd34479: data = 8'hfa;
      17'd34480: data = 8'hf6;
      17'd34481: data = 8'hf6;
      17'd34482: data = 8'hf9;
      17'd34483: data = 8'hfc;
      17'd34484: data = 8'hfe;
      17'd34485: data = 8'hfc;
      17'd34486: data = 8'hfc;
      17'd34487: data = 8'hfd;
      17'd34488: data = 8'h00;
      17'd34489: data = 8'h02;
      17'd34490: data = 8'h00;
      17'd34491: data = 8'h01;
      17'd34492: data = 8'h00;
      17'd34493: data = 8'hfe;
      17'd34494: data = 8'h06;
      17'd34495: data = 8'h05;
      17'd34496: data = 8'hfd;
      17'd34497: data = 8'h00;
      17'd34498: data = 8'hfd;
      17'd34499: data = 8'hfd;
      17'd34500: data = 8'h02;
      17'd34501: data = 8'hfd;
      17'd34502: data = 8'hfa;
      17'd34503: data = 8'h02;
      17'd34504: data = 8'hfd;
      17'd34505: data = 8'h11;
      17'd34506: data = 8'h0c;
      17'd34507: data = 8'hf5;
      17'd34508: data = 8'h0d;
      17'd34509: data = 8'h06;
      17'd34510: data = 8'h1a;
      17'd34511: data = 8'h15;
      17'd34512: data = 8'hf5;
      17'd34513: data = 8'h0a;
      17'd34514: data = 8'h0e;
      17'd34515: data = 8'h05;
      17'd34516: data = 8'hfe;
      17'd34517: data = 8'hf6;
      17'd34518: data = 8'h05;
      17'd34519: data = 8'hf6;
      17'd34520: data = 8'hfa;
      17'd34521: data = 8'h1a;
      17'd34522: data = 8'h04;
      17'd34523: data = 8'hf2;
      17'd34524: data = 8'h05;
      17'd34525: data = 8'h0d;
      17'd34526: data = 8'hfa;
      17'd34527: data = 8'h00;
      17'd34528: data = 8'h09;
      17'd34529: data = 8'hfa;
      17'd34530: data = 8'h05;
      17'd34531: data = 8'h09;
      17'd34532: data = 8'h05;
      17'd34533: data = 8'h00;
      17'd34534: data = 8'h04;
      17'd34535: data = 8'h01;
      17'd34536: data = 8'he9;
      17'd34537: data = 8'hfd;
      17'd34538: data = 8'h02;
      17'd34539: data = 8'hf2;
      17'd34540: data = 8'hfc;
      17'd34541: data = 8'h05;
      17'd34542: data = 8'h00;
      17'd34543: data = 8'hf9;
      17'd34544: data = 8'h0d;
      17'd34545: data = 8'h0a;
      17'd34546: data = 8'hfc;
      17'd34547: data = 8'h12;
      17'd34548: data = 8'h1e;
      17'd34549: data = 8'h16;
      17'd34550: data = 8'h16;
      17'd34551: data = 8'h13;
      17'd34552: data = 8'h1b;
      17'd34553: data = 8'h22;
      17'd34554: data = 8'h06;
      17'd34555: data = 8'h0e;
      17'd34556: data = 8'h04;
      17'd34557: data = 8'h05;
      17'd34558: data = 8'h0d;
      17'd34559: data = 8'hf5;
      17'd34560: data = 8'h02;
      17'd34561: data = 8'h09;
      17'd34562: data = 8'hf6;
      17'd34563: data = 8'hef;
      17'd34564: data = 8'hfe;
      17'd34565: data = 8'h01;
      17'd34566: data = 8'hf5;
      17'd34567: data = 8'hf5;
      17'd34568: data = 8'h04;
      17'd34569: data = 8'h02;
      17'd34570: data = 8'hfc;
      17'd34571: data = 8'h05;
      17'd34572: data = 8'hfe;
      17'd34573: data = 8'hf4;
      17'd34574: data = 8'hf4;
      17'd34575: data = 8'hf9;
      17'd34576: data = 8'hfa;
      17'd34577: data = 8'hfc;
      17'd34578: data = 8'hfa;
      17'd34579: data = 8'hf2;
      17'd34580: data = 8'h01;
      17'd34581: data = 8'h05;
      17'd34582: data = 8'hfd;
      17'd34583: data = 8'hfa;
      17'd34584: data = 8'hf6;
      17'd34585: data = 8'hfe;
      17'd34586: data = 8'h02;
      17'd34587: data = 8'h01;
      17'd34588: data = 8'h05;
      17'd34589: data = 8'h00;
      17'd34590: data = 8'hfe;
      17'd34591: data = 8'h02;
      17'd34592: data = 8'h01;
      17'd34593: data = 8'h00;
      17'd34594: data = 8'hfd;
      17'd34595: data = 8'hf4;
      17'd34596: data = 8'hfe;
      17'd34597: data = 8'h0a;
      17'd34598: data = 8'h00;
      17'd34599: data = 8'hfa;
      17'd34600: data = 8'h09;
      17'd34601: data = 8'h09;
      17'd34602: data = 8'hfd;
      17'd34603: data = 8'h04;
      17'd34604: data = 8'h0d;
      17'd34605: data = 8'h06;
      17'd34606: data = 8'h02;
      17'd34607: data = 8'h0d;
      17'd34608: data = 8'h15;
      17'd34609: data = 8'h06;
      17'd34610: data = 8'h0a;
      17'd34611: data = 8'h0a;
      17'd34612: data = 8'h05;
      17'd34613: data = 8'h0c;
      17'd34614: data = 8'h06;
      17'd34615: data = 8'h06;
      17'd34616: data = 8'h0c;
      17'd34617: data = 8'h0d;
      17'd34618: data = 8'h05;
      17'd34619: data = 8'h01;
      17'd34620: data = 8'h11;
      17'd34621: data = 8'h0c;
      17'd34622: data = 8'h00;
      17'd34623: data = 8'h09;
      17'd34624: data = 8'h0c;
      17'd34625: data = 8'h09;
      17'd34626: data = 8'h06;
      17'd34627: data = 8'h0a;
      17'd34628: data = 8'h0a;
      17'd34629: data = 8'h02;
      17'd34630: data = 8'h02;
      17'd34631: data = 8'h01;
      17'd34632: data = 8'h00;
      17'd34633: data = 8'hfd;
      17'd34634: data = 8'hf4;
      17'd34635: data = 8'hf4;
      17'd34636: data = 8'hfd;
      17'd34637: data = 8'hf9;
      17'd34638: data = 8'hf1;
      17'd34639: data = 8'hf5;
      17'd34640: data = 8'hfa;
      17'd34641: data = 8'hf6;
      17'd34642: data = 8'hf2;
      17'd34643: data = 8'hfa;
      17'd34644: data = 8'hfa;
      17'd34645: data = 8'hf5;
      17'd34646: data = 8'hfd;
      17'd34647: data = 8'h00;
      17'd34648: data = 8'hfe;
      17'd34649: data = 8'h00;
      17'd34650: data = 8'hfc;
      17'd34651: data = 8'hf9;
      17'd34652: data = 8'h00;
      17'd34653: data = 8'h01;
      17'd34654: data = 8'hfa;
      17'd34655: data = 8'hfc;
      17'd34656: data = 8'h00;
      17'd34657: data = 8'hfe;
      17'd34658: data = 8'hf9;
      17'd34659: data = 8'h00;
      17'd34660: data = 8'h00;
      17'd34661: data = 8'hed;
      17'd34662: data = 8'hef;
      17'd34663: data = 8'hfa;
      17'd34664: data = 8'hfc;
      17'd34665: data = 8'hf5;
      17'd34666: data = 8'hf4;
      17'd34667: data = 8'hf9;
      17'd34668: data = 8'hf2;
      17'd34669: data = 8'hed;
      17'd34670: data = 8'hf6;
      17'd34671: data = 8'hf2;
      17'd34672: data = 8'hed;
      17'd34673: data = 8'hef;
      17'd34674: data = 8'hf2;
      17'd34675: data = 8'hf6;
      17'd34676: data = 8'hf6;
      17'd34677: data = 8'he9;
      17'd34678: data = 8'heb;
      17'd34679: data = 8'hf6;
      17'd34680: data = 8'hf6;
      17'd34681: data = 8'hf2;
      17'd34682: data = 8'hf2;
      17'd34683: data = 8'hf5;
      17'd34684: data = 8'hfc;
      17'd34685: data = 8'hfd;
      17'd34686: data = 8'h02;
      17'd34687: data = 8'h05;
      17'd34688: data = 8'hf9;
      17'd34689: data = 8'hf5;
      17'd34690: data = 8'hf9;
      17'd34691: data = 8'hfc;
      17'd34692: data = 8'h00;
      17'd34693: data = 8'hf6;
      17'd34694: data = 8'hf1;
      17'd34695: data = 8'hfd;
      17'd34696: data = 8'hfa;
      17'd34697: data = 8'hf4;
      17'd34698: data = 8'hf5;
      17'd34699: data = 8'hf2;
      17'd34700: data = 8'hf5;
      17'd34701: data = 8'hf4;
      17'd34702: data = 8'hf6;
      17'd34703: data = 8'hf9;
      17'd34704: data = 8'hf2;
      17'd34705: data = 8'hef;
      17'd34706: data = 8'hf4;
      17'd34707: data = 8'hfd;
      17'd34708: data = 8'hf5;
      17'd34709: data = 8'he5;
      17'd34710: data = 8'hf2;
      17'd34711: data = 8'h01;
      17'd34712: data = 8'hfe;
      17'd34713: data = 8'hfe;
      17'd34714: data = 8'hf6;
      17'd34715: data = 8'hf2;
      17'd34716: data = 8'h0c;
      17'd34717: data = 8'h0d;
      17'd34718: data = 8'hf6;
      17'd34719: data = 8'hfc;
      17'd34720: data = 8'hf9;
      17'd34721: data = 8'h0a;
      17'd34722: data = 8'h27;
      17'd34723: data = 8'hfa;
      17'd34724: data = 8'hf1;
      17'd34725: data = 8'h05;
      17'd34726: data = 8'h11;
      17'd34727: data = 8'h13;
      17'd34728: data = 8'h0e;
      17'd34729: data = 8'h11;
      17'd34730: data = 8'he4;
      17'd34731: data = 8'hfd;
      17'd34732: data = 8'h33;
      17'd34733: data = 8'h05;
      17'd34734: data = 8'hed;
      17'd34735: data = 8'hfe;
      17'd34736: data = 8'hf4;
      17'd34737: data = 8'hfe;
      17'd34738: data = 8'h16;
      17'd34739: data = 8'hec;
      17'd34740: data = 8'hf9;
      17'd34741: data = 8'h19;
      17'd34742: data = 8'hd2;
      17'd34743: data = 8'hf4;
      17'd34744: data = 8'h34;
      17'd34745: data = 8'h11;
      17'd34746: data = 8'hde;
      17'd34747: data = 8'he9;
      17'd34748: data = 8'h29;
      17'd34749: data = 8'h0c;
      17'd34750: data = 8'h09;
      17'd34751: data = 8'h0e;
      17'd34752: data = 8'h00;
      17'd34753: data = 8'h05;
      17'd34754: data = 8'h04;
      17'd34755: data = 8'h19;
      17'd34756: data = 8'hf6;
      17'd34757: data = 8'h15;
      17'd34758: data = 8'h1f;
      17'd34759: data = 8'hd6;
      17'd34760: data = 8'h06;
      17'd34761: data = 8'h0d;
      17'd34762: data = 8'he7;
      17'd34763: data = 8'h0a;
      17'd34764: data = 8'h05;
      17'd34765: data = 8'hf5;
      17'd34766: data = 8'he9;
      17'd34767: data = 8'hfc;
      17'd34768: data = 8'h0a;
      17'd34769: data = 8'h02;
      17'd34770: data = 8'h05;
      17'd34771: data = 8'hde;
      17'd34772: data = 8'hf9;
      17'd34773: data = 8'h1a;
      17'd34774: data = 8'h09;
      17'd34775: data = 8'h15;
      17'd34776: data = 8'hfc;
      17'd34777: data = 8'hed;
      17'd34778: data = 8'h19;
      17'd34779: data = 8'h1a;
      17'd34780: data = 8'h04;
      17'd34781: data = 8'h19;
      17'd34782: data = 8'h05;
      17'd34783: data = 8'he9;
      17'd34784: data = 8'h0a;
      17'd34785: data = 8'h1f;
      17'd34786: data = 8'h13;
      17'd34787: data = 8'h0c;
      17'd34788: data = 8'hed;
      17'd34789: data = 8'hed;
      17'd34790: data = 8'h1b;
      17'd34791: data = 8'h1b;
      17'd34792: data = 8'h04;
      17'd34793: data = 8'h13;
      17'd34794: data = 8'h0c;
      17'd34795: data = 8'hf2;
      17'd34796: data = 8'h09;
      17'd34797: data = 8'h16;
      17'd34798: data = 8'h05;
      17'd34799: data = 8'h00;
      17'd34800: data = 8'hf9;
      17'd34801: data = 8'h01;
      17'd34802: data = 8'h0e;
      17'd34803: data = 8'hfa;
      17'd34804: data = 8'h00;
      17'd34805: data = 8'h0e;
      17'd34806: data = 8'hef;
      17'd34807: data = 8'hec;
      17'd34808: data = 8'h04;
      17'd34809: data = 8'hfe;
      17'd34810: data = 8'h0d;
      17'd34811: data = 8'h0d;
      17'd34812: data = 8'hf1;
      17'd34813: data = 8'hf9;
      17'd34814: data = 8'h13;
      17'd34815: data = 8'h1b;
      17'd34816: data = 8'h0e;
      17'd34817: data = 8'h00;
      17'd34818: data = 8'hfe;
      17'd34819: data = 8'h05;
      17'd34820: data = 8'h13;
      17'd34821: data = 8'h19;
      17'd34822: data = 8'h12;
      17'd34823: data = 8'hfe;
      17'd34824: data = 8'hed;
      17'd34825: data = 8'h01;
      17'd34826: data = 8'h13;
      17'd34827: data = 8'h01;
      17'd34828: data = 8'hf4;
      17'd34829: data = 8'hfc;
      17'd34830: data = 8'hf5;
      17'd34831: data = 8'hfd;
      17'd34832: data = 8'h12;
      17'd34833: data = 8'h06;
      17'd34834: data = 8'hf1;
      17'd34835: data = 8'hf4;
      17'd34836: data = 8'h02;
      17'd34837: data = 8'h11;
      17'd34838: data = 8'h0a;
      17'd34839: data = 8'h01;
      17'd34840: data = 8'hfd;
      17'd34841: data = 8'hf6;
      17'd34842: data = 8'h02;
      17'd34843: data = 8'h09;
      17'd34844: data = 8'hfd;
      17'd34845: data = 8'hfe;
      17'd34846: data = 8'hf5;
      17'd34847: data = 8'hf2;
      17'd34848: data = 8'h05;
      17'd34849: data = 8'h0d;
      17'd34850: data = 8'hf9;
      17'd34851: data = 8'hf2;
      17'd34852: data = 8'h0d;
      17'd34853: data = 8'h09;
      17'd34854: data = 8'hfd;
      17'd34855: data = 8'hfe;
      17'd34856: data = 8'h02;
      17'd34857: data = 8'h04;
      17'd34858: data = 8'h09;
      17'd34859: data = 8'h0e;
      17'd34860: data = 8'h00;
      17'd34861: data = 8'hef;
      17'd34862: data = 8'h02;
      17'd34863: data = 8'h0e;
      17'd34864: data = 8'hf6;
      17'd34865: data = 8'hf5;
      17'd34866: data = 8'hfa;
      17'd34867: data = 8'hfe;
      17'd34868: data = 8'h12;
      17'd34869: data = 8'hfd;
      17'd34870: data = 8'he4;
      17'd34871: data = 8'hfa;
      17'd34872: data = 8'h02;
      17'd34873: data = 8'hfc;
      17'd34874: data = 8'hfe;
      17'd34875: data = 8'hfd;
      17'd34876: data = 8'he7;
      17'd34877: data = 8'hf2;
      17'd34878: data = 8'h04;
      17'd34879: data = 8'h02;
      17'd34880: data = 8'hfd;
      17'd34881: data = 8'hf2;
      17'd34882: data = 8'hec;
      17'd34883: data = 8'hfa;
      17'd34884: data = 8'h13;
      17'd34885: data = 8'hfe;
      17'd34886: data = 8'he0;
      17'd34887: data = 8'h00;
      17'd34888: data = 8'h19;
      17'd34889: data = 8'h00;
      17'd34890: data = 8'hfa;
      17'd34891: data = 8'h04;
      17'd34892: data = 8'hfa;
      17'd34893: data = 8'hfc;
      17'd34894: data = 8'h04;
      17'd34895: data = 8'hf6;
      17'd34896: data = 8'hf6;
      17'd34897: data = 8'h11;
      17'd34898: data = 8'hf2;
      17'd34899: data = 8'hd8;
      17'd34900: data = 8'h06;
      17'd34901: data = 8'h00;
      17'd34902: data = 8'he9;
      17'd34903: data = 8'h02;
      17'd34904: data = 8'heb;
      17'd34905: data = 8'he0;
      17'd34906: data = 8'h02;
      17'd34907: data = 8'h00;
      17'd34908: data = 8'hfa;
      17'd34909: data = 8'h02;
      17'd34910: data = 8'he5;
      17'd34911: data = 8'he0;
      17'd34912: data = 8'h06;
      17'd34913: data = 8'h22;
      17'd34914: data = 8'h06;
      17'd34915: data = 8'hd5;
      17'd34916: data = 8'he9;
      17'd34917: data = 8'h1b;
      17'd34918: data = 8'h0e;
      17'd34919: data = 8'hfd;
      17'd34920: data = 8'h02;
      17'd34921: data = 8'hec;
      17'd34922: data = 8'hfc;
      17'd34923: data = 8'h05;
      17'd34924: data = 8'hfa;
      17'd34925: data = 8'h23;
      17'd34926: data = 8'hfa;
      17'd34927: data = 8'hce;
      17'd34928: data = 8'h0d;
      17'd34929: data = 8'h0d;
      17'd34930: data = 8'hec;
      17'd34931: data = 8'h09;
      17'd34932: data = 8'h00;
      17'd34933: data = 8'hd8;
      17'd34934: data = 8'hf6;
      17'd34935: data = 8'h16;
      17'd34936: data = 8'he9;
      17'd34937: data = 8'hf2;
      17'd34938: data = 8'hfd;
      17'd34939: data = 8'hde;
      17'd34940: data = 8'h15;
      17'd34941: data = 8'h05;
      17'd34942: data = 8'hd6;
      17'd34943: data = 8'hfa;
      17'd34944: data = 8'h19;
      17'd34945: data = 8'hf5;
      17'd34946: data = 8'hf2;
      17'd34947: data = 8'h11;
      17'd34948: data = 8'hf2;
      17'd34949: data = 8'hf6;
      17'd34950: data = 8'hf1;
      17'd34951: data = 8'hf1;
      17'd34952: data = 8'h1b;
      17'd34953: data = 8'h01;
      17'd34954: data = 8'hd8;
      17'd34955: data = 8'hfe;
      17'd34956: data = 8'h1b;
      17'd34957: data = 8'hf1;
      17'd34958: data = 8'hfd;
      17'd34959: data = 8'h04;
      17'd34960: data = 8'hed;
      17'd34961: data = 8'h00;
      17'd34962: data = 8'h1f;
      17'd34963: data = 8'h05;
      17'd34964: data = 8'hd1;
      17'd34965: data = 8'h02;
      17'd34966: data = 8'h24;
      17'd34967: data = 8'hdc;
      17'd34968: data = 8'h02;
      17'd34969: data = 8'h33;
      17'd34970: data = 8'hbd;
      17'd34971: data = 8'hef;
      17'd34972: data = 8'h1e;
      17'd34973: data = 8'hca;
      17'd34974: data = 8'h1e;
      17'd34975: data = 8'h12;
      17'd34976: data = 8'hc5;
      17'd34977: data = 8'h0e;
      17'd34978: data = 8'h04;
      17'd34979: data = 8'hef;
      17'd34980: data = 8'h06;
      17'd34981: data = 8'h09;
      17'd34982: data = 8'h1a;
      17'd34983: data = 8'hf1;
      17'd34984: data = 8'he0;
      17'd34985: data = 8'h23;
      17'd34986: data = 8'h0c;
      17'd34987: data = 8'hef;
      17'd34988: data = 8'h13;
      17'd34989: data = 8'hfc;
      17'd34990: data = 8'hf1;
      17'd34991: data = 8'h1a;
      17'd34992: data = 8'hf9;
      17'd34993: data = 8'hec;
      17'd34994: data = 8'h11;
      17'd34995: data = 8'h02;
      17'd34996: data = 8'hf9;
      17'd34997: data = 8'h00;
      17'd34998: data = 8'hec;
      17'd34999: data = 8'hf4;
      17'd35000: data = 8'h1f;
      17'd35001: data = 8'hfc;
      17'd35002: data = 8'he7;
      17'd35003: data = 8'h09;
      17'd35004: data = 8'he9;
      17'd35005: data = 8'h02;
      17'd35006: data = 8'h24;
      17'd35007: data = 8'hde;
      17'd35008: data = 8'hef;
      17'd35009: data = 8'h12;
      17'd35010: data = 8'hfc;
      17'd35011: data = 8'h16;
      17'd35012: data = 8'h01;
      17'd35013: data = 8'hec;
      17'd35014: data = 8'h12;
      17'd35015: data = 8'h01;
      17'd35016: data = 8'h05;
      17'd35017: data = 8'h23;
      17'd35018: data = 8'h04;
      17'd35019: data = 8'hfa;
      17'd35020: data = 8'h01;
      17'd35021: data = 8'h0d;
      17'd35022: data = 8'h23;
      17'd35023: data = 8'h05;
      17'd35024: data = 8'h04;
      17'd35025: data = 8'h06;
      17'd35026: data = 8'hf2;
      17'd35027: data = 8'h09;
      17'd35028: data = 8'h11;
      17'd35029: data = 8'h1a;
      17'd35030: data = 8'h04;
      17'd35031: data = 8'hd3;
      17'd35032: data = 8'h02;
      17'd35033: data = 8'h31;
      17'd35034: data = 8'hfe;
      17'd35035: data = 8'hf1;
      17'd35036: data = 8'hfa;
      17'd35037: data = 8'hfe;
      17'd35038: data = 8'h16;
      17'd35039: data = 8'h26;
      17'd35040: data = 8'he9;
      17'd35041: data = 8'hd5;
      17'd35042: data = 8'h2b;
      17'd35043: data = 8'h09;
      17'd35044: data = 8'hf4;
      17'd35045: data = 8'h23;
      17'd35046: data = 8'hf2;
      17'd35047: data = 8'hfe;
      17'd35048: data = 8'h1b;
      17'd35049: data = 8'hf5;
      17'd35050: data = 8'h0c;
      17'd35051: data = 8'h15;
      17'd35052: data = 8'hf9;
      17'd35053: data = 8'h15;
      17'd35054: data = 8'h1a;
      17'd35055: data = 8'hf6;
      17'd35056: data = 8'h05;
      17'd35057: data = 8'h13;
      17'd35058: data = 8'h1a;
      17'd35059: data = 8'hf6;
      17'd35060: data = 8'hf4;
      17'd35061: data = 8'h0c;
      17'd35062: data = 8'h02;
      17'd35063: data = 8'h09;
      17'd35064: data = 8'hfa;
      17'd35065: data = 8'hef;
      17'd35066: data = 8'hfe;
      17'd35067: data = 8'h04;
      17'd35068: data = 8'h04;
      17'd35069: data = 8'hfc;
      17'd35070: data = 8'hf5;
      17'd35071: data = 8'hfa;
      17'd35072: data = 8'h05;
      17'd35073: data = 8'h04;
      17'd35074: data = 8'hfd;
      17'd35075: data = 8'h04;
      17'd35076: data = 8'hf5;
      17'd35077: data = 8'h00;
      17'd35078: data = 8'h16;
      17'd35079: data = 8'h00;
      17'd35080: data = 8'hf4;
      17'd35081: data = 8'h09;
      17'd35082: data = 8'h0c;
      17'd35083: data = 8'hfa;
      17'd35084: data = 8'h00;
      17'd35085: data = 8'h09;
      17'd35086: data = 8'h0c;
      17'd35087: data = 8'h04;
      17'd35088: data = 8'hf6;
      17'd35089: data = 8'h00;
      17'd35090: data = 8'h00;
      17'd35091: data = 8'h00;
      17'd35092: data = 8'h1b;
      17'd35093: data = 8'hfc;
      17'd35094: data = 8'he3;
      17'd35095: data = 8'h11;
      17'd35096: data = 8'h04;
      17'd35097: data = 8'hf4;
      17'd35098: data = 8'hfc;
      17'd35099: data = 8'heb;
      17'd35100: data = 8'hfe;
      17'd35101: data = 8'h04;
      17'd35102: data = 8'hf2;
      17'd35103: data = 8'hf1;
      17'd35104: data = 8'hfd;
      17'd35105: data = 8'hf6;
      17'd35106: data = 8'hf6;
      17'd35107: data = 8'h09;
      17'd35108: data = 8'hef;
      17'd35109: data = 8'hde;
      17'd35110: data = 8'hfe;
      17'd35111: data = 8'h0d;
      17'd35112: data = 8'he5;
      17'd35113: data = 8'hed;
      17'd35114: data = 8'h12;
      17'd35115: data = 8'hf5;
      17'd35116: data = 8'heb;
      17'd35117: data = 8'h0d;
      17'd35118: data = 8'hfc;
      17'd35119: data = 8'he4;
      17'd35120: data = 8'h0d;
      17'd35121: data = 8'h0d;
      17'd35122: data = 8'hef;
      17'd35123: data = 8'h04;
      17'd35124: data = 8'h04;
      17'd35125: data = 8'hef;
      17'd35126: data = 8'hfd;
      17'd35127: data = 8'h0c;
      17'd35128: data = 8'hf5;
      17'd35129: data = 8'he5;
      17'd35130: data = 8'hfe;
      17'd35131: data = 8'hfe;
      17'd35132: data = 8'hf4;
      17'd35133: data = 8'hfe;
      17'd35134: data = 8'hf9;
      17'd35135: data = 8'he7;
      17'd35136: data = 8'hf6;
      17'd35137: data = 8'hfe;
      17'd35138: data = 8'hf5;
      17'd35139: data = 8'hf9;
      17'd35140: data = 8'hf4;
      17'd35141: data = 8'he4;
      17'd35142: data = 8'hfc;
      17'd35143: data = 8'h15;
      17'd35144: data = 8'hf6;
      17'd35145: data = 8'he3;
      17'd35146: data = 8'hf6;
      17'd35147: data = 8'h00;
      17'd35148: data = 8'h00;
      17'd35149: data = 8'h02;
      17'd35150: data = 8'h04;
      17'd35151: data = 8'hef;
      17'd35152: data = 8'hf5;
      17'd35153: data = 8'h19;
      17'd35154: data = 8'h02;
      17'd35155: data = 8'he9;
      17'd35156: data = 8'hfe;
      17'd35157: data = 8'h06;
      17'd35158: data = 8'hfd;
      17'd35159: data = 8'hf1;
      17'd35160: data = 8'hf4;
      17'd35161: data = 8'hfe;
      17'd35162: data = 8'h05;
      17'd35163: data = 8'h00;
      17'd35164: data = 8'he9;
      17'd35165: data = 8'hec;
      17'd35166: data = 8'h06;
      17'd35167: data = 8'h06;
      17'd35168: data = 8'he3;
      17'd35169: data = 8'hf9;
      17'd35170: data = 8'h0e;
      17'd35171: data = 8'he9;
      17'd35172: data = 8'hfa;
      17'd35173: data = 8'h0d;
      17'd35174: data = 8'he0;
      17'd35175: data = 8'hf6;
      17'd35176: data = 8'h13;
      17'd35177: data = 8'he9;
      17'd35178: data = 8'h0a;
      17'd35179: data = 8'h04;
      17'd35180: data = 8'he0;
      17'd35181: data = 8'h1f;
      17'd35182: data = 8'h0d;
      17'd35183: data = 8'hd5;
      17'd35184: data = 8'hf5;
      17'd35185: data = 8'h2b;
      17'd35186: data = 8'h04;
      17'd35187: data = 8'hd6;
      17'd35188: data = 8'h00;
      17'd35189: data = 8'hf9;
      17'd35190: data = 8'h09;
      17'd35191: data = 8'h23;
      17'd35192: data = 8'he3;
      17'd35193: data = 8'hd8;
      17'd35194: data = 8'h0a;
      17'd35195: data = 8'h12;
      17'd35196: data = 8'h0d;
      17'd35197: data = 8'hf4;
      17'd35198: data = 8'hd6;
      17'd35199: data = 8'h0d;
      17'd35200: data = 8'h2b;
      17'd35201: data = 8'hf2;
      17'd35202: data = 8'he5;
      17'd35203: data = 8'h04;
      17'd35204: data = 8'h02;
      17'd35205: data = 8'hf5;
      17'd35206: data = 8'hfe;
      17'd35207: data = 8'h06;
      17'd35208: data = 8'hef;
      17'd35209: data = 8'h02;
      17'd35210: data = 8'h0c;
      17'd35211: data = 8'hed;
      17'd35212: data = 8'h04;
      17'd35213: data = 8'h00;
      17'd35214: data = 8'h04;
      17'd35215: data = 8'h1e;
      17'd35216: data = 8'hed;
      17'd35217: data = 8'hec;
      17'd35218: data = 8'h19;
      17'd35219: data = 8'h15;
      17'd35220: data = 8'hfa;
      17'd35221: data = 8'hef;
      17'd35222: data = 8'hfa;
      17'd35223: data = 8'h0e;
      17'd35224: data = 8'h12;
      17'd35225: data = 8'he9;
      17'd35226: data = 8'hfc;
      17'd35227: data = 8'h00;
      17'd35228: data = 8'hf9;
      17'd35229: data = 8'h0d;
      17'd35230: data = 8'hf1;
      17'd35231: data = 8'h0e;
      17'd35232: data = 8'h0e;
      17'd35233: data = 8'hcd;
      17'd35234: data = 8'h06;
      17'd35235: data = 8'h22;
      17'd35236: data = 8'hf5;
      17'd35237: data = 8'h0a;
      17'd35238: data = 8'hf5;
      17'd35239: data = 8'hde;
      17'd35240: data = 8'h0a;
      17'd35241: data = 8'h23;
      17'd35242: data = 8'h06;
      17'd35243: data = 8'hcd;
      17'd35244: data = 8'hdc;
      17'd35245: data = 8'h34;
      17'd35246: data = 8'h22;
      17'd35247: data = 8'hc6;
      17'd35248: data = 8'hfc;
      17'd35249: data = 8'h11;
      17'd35250: data = 8'hdc;
      17'd35251: data = 8'h24;
      17'd35252: data = 8'h2f;
      17'd35253: data = 8'hd2;
      17'd35254: data = 8'hdc;
      17'd35255: data = 8'h31;
      17'd35256: data = 8'h16;
      17'd35257: data = 8'hef;
      17'd35258: data = 8'h0a;
      17'd35259: data = 8'h12;
      17'd35260: data = 8'hf6;
      17'd35261: data = 8'hfa;
      17'd35262: data = 8'h2f;
      17'd35263: data = 8'hec;
      17'd35264: data = 8'hc9;
      17'd35265: data = 8'h34;
      17'd35266: data = 8'h19;
      17'd35267: data = 8'hed;
      17'd35268: data = 8'he4;
      17'd35269: data = 8'hf9;
      17'd35270: data = 8'h34;
      17'd35271: data = 8'hf1;
      17'd35272: data = 8'he2;
      17'd35273: data = 8'h1a;
      17'd35274: data = 8'h02;
      17'd35275: data = 8'hf5;
      17'd35276: data = 8'hfd;
      17'd35277: data = 8'hfd;
      17'd35278: data = 8'h0e;
      17'd35279: data = 8'h02;
      17'd35280: data = 8'h16;
      17'd35281: data = 8'hfa;
      17'd35282: data = 8'hcd;
      17'd35283: data = 8'h1f;
      17'd35284: data = 8'h2f;
      17'd35285: data = 8'h11;
      17'd35286: data = 8'he2;
      17'd35287: data = 8'he0;
      17'd35288: data = 8'h24;
      17'd35289: data = 8'h2d;
      17'd35290: data = 8'h11;
      17'd35291: data = 8'hd5;
      17'd35292: data = 8'hf4;
      17'd35293: data = 8'h26;
      17'd35294: data = 8'h13;
      17'd35295: data = 8'h05;
      17'd35296: data = 8'heb;
      17'd35297: data = 8'hde;
      17'd35298: data = 8'h15;
      17'd35299: data = 8'h43;
      17'd35300: data = 8'he0;
      17'd35301: data = 8'hbc;
      17'd35302: data = 8'h12;
      17'd35303: data = 8'h1c;
      17'd35304: data = 8'h13;
      17'd35305: data = 8'hed;
      17'd35306: data = 8'hdc;
      17'd35307: data = 8'h0a;
      17'd35308: data = 8'h0e;
      17'd35309: data = 8'h05;
      17'd35310: data = 8'hfc;
      17'd35311: data = 8'hef;
      17'd35312: data = 8'h0d;
      17'd35313: data = 8'h05;
      17'd35314: data = 8'hfc;
      17'd35315: data = 8'h06;
      17'd35316: data = 8'hf1;
      17'd35317: data = 8'h05;
      17'd35318: data = 8'h22;
      17'd35319: data = 8'h00;
      17'd35320: data = 8'hde;
      17'd35321: data = 8'h02;
      17'd35322: data = 8'h1a;
      17'd35323: data = 8'hf5;
      17'd35324: data = 8'h16;
      17'd35325: data = 8'h05;
      17'd35326: data = 8'hd5;
      17'd35327: data = 8'h1b;
      17'd35328: data = 8'h2f;
      17'd35329: data = 8'he3;
      17'd35330: data = 8'he3;
      17'd35331: data = 8'h0d;
      17'd35332: data = 8'h1f;
      17'd35333: data = 8'h09;
      17'd35334: data = 8'hdb;
      17'd35335: data = 8'hf9;
      17'd35336: data = 8'h13;
      17'd35337: data = 8'hfd;
      17'd35338: data = 8'h02;
      17'd35339: data = 8'h11;
      17'd35340: data = 8'hde;
      17'd35341: data = 8'hec;
      17'd35342: data = 8'h2d;
      17'd35343: data = 8'hfe;
      17'd35344: data = 8'hd2;
      17'd35345: data = 8'h05;
      17'd35346: data = 8'h05;
      17'd35347: data = 8'h13;
      17'd35348: data = 8'h0c;
      17'd35349: data = 8'hbc;
      17'd35350: data = 8'hf4;
      17'd35351: data = 8'h3a;
      17'd35352: data = 8'hec;
      17'd35353: data = 8'he5;
      17'd35354: data = 8'h19;
      17'd35355: data = 8'he2;
      17'd35356: data = 8'heb;
      17'd35357: data = 8'h35;
      17'd35358: data = 8'h02;
      17'd35359: data = 8'hce;
      17'd35360: data = 8'h0d;
      17'd35361: data = 8'h1a;
      17'd35362: data = 8'h02;
      17'd35363: data = 8'hf6;
      17'd35364: data = 8'he5;
      17'd35365: data = 8'h11;
      17'd35366: data = 8'h1c;
      17'd35367: data = 8'heb;
      17'd35368: data = 8'he9;
      17'd35369: data = 8'h16;
      17'd35370: data = 8'hf5;
      17'd35371: data = 8'hd5;
      17'd35372: data = 8'h13;
      17'd35373: data = 8'h23;
      17'd35374: data = 8'hdc;
      17'd35375: data = 8'he9;
      17'd35376: data = 8'h0a;
      17'd35377: data = 8'hfa;
      17'd35378: data = 8'h05;
      17'd35379: data = 8'hfe;
      17'd35380: data = 8'he9;
      17'd35381: data = 8'h02;
      17'd35382: data = 8'h05;
      17'd35383: data = 8'hfd;
      17'd35384: data = 8'hfd;
      17'd35385: data = 8'hec;
      17'd35386: data = 8'h02;
      17'd35387: data = 8'h01;
      17'd35388: data = 8'he9;
      17'd35389: data = 8'h19;
      17'd35390: data = 8'h09;
      17'd35391: data = 8'hc2;
      17'd35392: data = 8'h0d;
      17'd35393: data = 8'h1a;
      17'd35394: data = 8'hec;
      17'd35395: data = 8'h0d;
      17'd35396: data = 8'hf5;
      17'd35397: data = 8'he2;
      17'd35398: data = 8'h1e;
      17'd35399: data = 8'h09;
      17'd35400: data = 8'he2;
      17'd35401: data = 8'hfc;
      17'd35402: data = 8'h04;
      17'd35403: data = 8'h19;
      17'd35404: data = 8'h04;
      17'd35405: data = 8'hda;
      17'd35406: data = 8'hf2;
      17'd35407: data = 8'h05;
      17'd35408: data = 8'h05;
      17'd35409: data = 8'h0c;
      17'd35410: data = 8'hed;
      17'd35411: data = 8'hd1;
      17'd35412: data = 8'h09;
      17'd35413: data = 8'h1a;
      17'd35414: data = 8'he5;
      17'd35415: data = 8'h09;
      17'd35416: data = 8'hf6;
      17'd35417: data = 8'hde;
      17'd35418: data = 8'h23;
      17'd35419: data = 8'h15;
      17'd35420: data = 8'hd6;
      17'd35421: data = 8'hf6;
      17'd35422: data = 8'h16;
      17'd35423: data = 8'h01;
      17'd35424: data = 8'hfe;
      17'd35425: data = 8'hf1;
      17'd35426: data = 8'hed;
      17'd35427: data = 8'h0d;
      17'd35428: data = 8'hfd;
      17'd35429: data = 8'hfc;
      17'd35430: data = 8'hfa;
      17'd35431: data = 8'heb;
      17'd35432: data = 8'h05;
      17'd35433: data = 8'h0e;
      17'd35434: data = 8'hf9;
      17'd35435: data = 8'h04;
      17'd35436: data = 8'hf2;
      17'd35437: data = 8'he5;
      17'd35438: data = 8'h27;
      17'd35439: data = 8'h0e;
      17'd35440: data = 8'hda;
      17'd35441: data = 8'he5;
      17'd35442: data = 8'h19;
      17'd35443: data = 8'h1a;
      17'd35444: data = 8'he0;
      17'd35445: data = 8'hf4;
      17'd35446: data = 8'hfd;
      17'd35447: data = 8'h04;
      17'd35448: data = 8'h09;
      17'd35449: data = 8'he2;
      17'd35450: data = 8'h0a;
      17'd35451: data = 8'h0d;
      17'd35452: data = 8'he4;
      17'd35453: data = 8'h04;
      17'd35454: data = 8'h26;
      17'd35455: data = 8'heb;
      17'd35456: data = 8'hc9;
      17'd35457: data = 8'h1c;
      17'd35458: data = 8'h1e;
      17'd35459: data = 8'hf1;
      17'd35460: data = 8'he7;
      17'd35461: data = 8'hf5;
      17'd35462: data = 8'h00;
      17'd35463: data = 8'h13;
      17'd35464: data = 8'h0c;
      17'd35465: data = 8'hd6;
      17'd35466: data = 8'h05;
      17'd35467: data = 8'h19;
      17'd35468: data = 8'hf2;
      17'd35469: data = 8'hfa;
      17'd35470: data = 8'h00;
      17'd35471: data = 8'hfc;
      17'd35472: data = 8'h0c;
      17'd35473: data = 8'h06;
      17'd35474: data = 8'hed;
      17'd35475: data = 8'hfe;
      17'd35476: data = 8'hef;
      17'd35477: data = 8'h00;
      17'd35478: data = 8'h1c;
      17'd35479: data = 8'hfe;
      17'd35480: data = 8'he3;
      17'd35481: data = 8'heb;
      17'd35482: data = 8'h0d;
      17'd35483: data = 8'h0d;
      17'd35484: data = 8'he9;
      17'd35485: data = 8'he9;
      17'd35486: data = 8'h15;
      17'd35487: data = 8'hfe;
      17'd35488: data = 8'hde;
      17'd35489: data = 8'h00;
      17'd35490: data = 8'h0d;
      17'd35491: data = 8'hfd;
      17'd35492: data = 8'h0d;
      17'd35493: data = 8'hf5;
      17'd35494: data = 8'hec;
      17'd35495: data = 8'h19;
      17'd35496: data = 8'h05;
      17'd35497: data = 8'h0c;
      17'd35498: data = 8'h11;
      17'd35499: data = 8'heb;
      17'd35500: data = 8'hfc;
      17'd35501: data = 8'h29;
      17'd35502: data = 8'h1a;
      17'd35503: data = 8'hdb;
      17'd35504: data = 8'hf9;
      17'd35505: data = 8'h1b;
      17'd35506: data = 8'h09;
      17'd35507: data = 8'h00;
      17'd35508: data = 8'h04;
      17'd35509: data = 8'hed;
      17'd35510: data = 8'hed;
      17'd35511: data = 8'h1a;
      17'd35512: data = 8'h04;
      17'd35513: data = 8'h00;
      17'd35514: data = 8'hf5;
      17'd35515: data = 8'hf5;
      17'd35516: data = 8'hf9;
      17'd35517: data = 8'h09;
      17'd35518: data = 8'h16;
      17'd35519: data = 8'hef;
      17'd35520: data = 8'h02;
      17'd35521: data = 8'h13;
      17'd35522: data = 8'heb;
      17'd35523: data = 8'h15;
      17'd35524: data = 8'h1a;
      17'd35525: data = 8'hf2;
      17'd35526: data = 8'h11;
      17'd35527: data = 8'h05;
      17'd35528: data = 8'h12;
      17'd35529: data = 8'hef;
      17'd35530: data = 8'h11;
      17'd35531: data = 8'h22;
      17'd35532: data = 8'he5;
      17'd35533: data = 8'h0d;
      17'd35534: data = 8'hed;
      17'd35535: data = 8'h00;
      17'd35536: data = 8'h2b;
      17'd35537: data = 8'hf9;
      17'd35538: data = 8'hef;
      17'd35539: data = 8'hed;
      17'd35540: data = 8'h11;
      17'd35541: data = 8'h06;
      17'd35542: data = 8'hfc;
      17'd35543: data = 8'h0c;
      17'd35544: data = 8'he9;
      17'd35545: data = 8'h09;
      17'd35546: data = 8'h0a;
      17'd35547: data = 8'hed;
      17'd35548: data = 8'h0d;
      17'd35549: data = 8'h06;
      17'd35550: data = 8'hfe;
      17'd35551: data = 8'h00;
      17'd35552: data = 8'h0a;
      17'd35553: data = 8'hfe;
      17'd35554: data = 8'hf9;
      17'd35555: data = 8'h1b;
      17'd35556: data = 8'h04;
      17'd35557: data = 8'hed;
      17'd35558: data = 8'h24;
      17'd35559: data = 8'hfc;
      17'd35560: data = 8'he5;
      17'd35561: data = 8'h3d;
      17'd35562: data = 8'h04;
      17'd35563: data = 8'hda;
      17'd35564: data = 8'h1a;
      17'd35565: data = 8'h12;
      17'd35566: data = 8'hfe;
      17'd35567: data = 8'h0a;
      17'd35568: data = 8'hef;
      17'd35569: data = 8'hfe;
      17'd35570: data = 8'h1a;
      17'd35571: data = 8'hf1;
      17'd35572: data = 8'hfa;
      17'd35573: data = 8'h0c;
      17'd35574: data = 8'hf6;
      17'd35575: data = 8'hf2;
      17'd35576: data = 8'h01;
      17'd35577: data = 8'h0a;
      17'd35578: data = 8'hf4;
      17'd35579: data = 8'hfe;
      17'd35580: data = 8'hf9;
      17'd35581: data = 8'hec;
      17'd35582: data = 8'h23;
      17'd35583: data = 8'h04;
      17'd35584: data = 8'hcb;
      17'd35585: data = 8'h11;
      17'd35586: data = 8'h16;
      17'd35587: data = 8'hfa;
      17'd35588: data = 8'hec;
      17'd35589: data = 8'hfd;
      17'd35590: data = 8'h12;
      17'd35591: data = 8'h02;
      17'd35592: data = 8'h01;
      17'd35593: data = 8'hf6;
      17'd35594: data = 8'hfd;
      17'd35595: data = 8'h16;
      17'd35596: data = 8'h1e;
      17'd35597: data = 8'hd6;
      17'd35598: data = 8'h01;
      17'd35599: data = 8'h23;
      17'd35600: data = 8'hf4;
      17'd35601: data = 8'h11;
      17'd35602: data = 8'h11;
      17'd35603: data = 8'he2;
      17'd35604: data = 8'hf5;
      17'd35605: data = 8'h1f;
      17'd35606: data = 8'h23;
      17'd35607: data = 8'heb;
      17'd35608: data = 8'hc9;
      17'd35609: data = 8'h0e;
      17'd35610: data = 8'h1e;
      17'd35611: data = 8'h01;
      17'd35612: data = 8'he7;
      17'd35613: data = 8'he3;
      17'd35614: data = 8'h1c;
      17'd35615: data = 8'h02;
      17'd35616: data = 8'he4;
      17'd35617: data = 8'h09;
      17'd35618: data = 8'he9;
      17'd35619: data = 8'hf1;
      17'd35620: data = 8'h35;
      17'd35621: data = 8'he5;
      17'd35622: data = 8'hd2;
      17'd35623: data = 8'h29;
      17'd35624: data = 8'hfa;
      17'd35625: data = 8'hfc;
      17'd35626: data = 8'h0a;
      17'd35627: data = 8'hec;
      17'd35628: data = 8'h06;
      17'd35629: data = 8'h1a;
      17'd35630: data = 8'hf5;
      17'd35631: data = 8'he7;
      17'd35632: data = 8'h15;
      17'd35633: data = 8'hfc;
      17'd35634: data = 8'hed;
      17'd35635: data = 8'h2d;
      17'd35636: data = 8'hfc;
      17'd35637: data = 8'hc2;
      17'd35638: data = 8'h13;
      17'd35639: data = 8'h24;
      17'd35640: data = 8'he2;
      17'd35641: data = 8'h05;
      17'd35642: data = 8'h16;
      17'd35643: data = 8'hd1;
      17'd35644: data = 8'hfe;
      17'd35645: data = 8'h24;
      17'd35646: data = 8'heb;
      17'd35647: data = 8'hef;
      17'd35648: data = 8'h16;
      17'd35649: data = 8'heb;
      17'd35650: data = 8'he3;
      17'd35651: data = 8'h05;
      17'd35652: data = 8'h12;
      17'd35653: data = 8'h0a;
      17'd35654: data = 8'hda;
      17'd35655: data = 8'hde;
      17'd35656: data = 8'h19;
      17'd35657: data = 8'h22;
      17'd35658: data = 8'hf5;
      17'd35659: data = 8'heb;
      17'd35660: data = 8'hf6;
      17'd35661: data = 8'h0c;
      17'd35662: data = 8'h16;
      17'd35663: data = 8'hfc;
      17'd35664: data = 8'hf5;
      17'd35665: data = 8'hfc;
      17'd35666: data = 8'hfe;
      17'd35667: data = 8'h19;
      17'd35668: data = 8'h05;
      17'd35669: data = 8'heb;
      17'd35670: data = 8'h04;
      17'd35671: data = 8'hf5;
      17'd35672: data = 8'hf6;
      17'd35673: data = 8'h23;
      17'd35674: data = 8'hf4;
      17'd35675: data = 8'he2;
      17'd35676: data = 8'h00;
      17'd35677: data = 8'h05;
      17'd35678: data = 8'h04;
      17'd35679: data = 8'h01;
      17'd35680: data = 8'hf5;
      17'd35681: data = 8'hfe;
      17'd35682: data = 8'hf1;
      17'd35683: data = 8'h15;
      17'd35684: data = 8'h09;
      17'd35685: data = 8'hd2;
      17'd35686: data = 8'h1a;
      17'd35687: data = 8'h0c;
      17'd35688: data = 8'hf1;
      17'd35689: data = 8'h11;
      17'd35690: data = 8'hed;
      17'd35691: data = 8'hde;
      17'd35692: data = 8'h0e;
      17'd35693: data = 8'h05;
      17'd35694: data = 8'hfc;
      17'd35695: data = 8'hec;
      17'd35696: data = 8'he3;
      17'd35697: data = 8'h00;
      17'd35698: data = 8'h01;
      17'd35699: data = 8'h0c;
      17'd35700: data = 8'hfe;
      17'd35701: data = 8'he2;
      17'd35702: data = 8'hf6;
      17'd35703: data = 8'h13;
      17'd35704: data = 8'h06;
      17'd35705: data = 8'hf1;
      17'd35706: data = 8'h04;
      17'd35707: data = 8'h0d;
      17'd35708: data = 8'he2;
      17'd35709: data = 8'h0e;
      17'd35710: data = 8'h16;
      17'd35711: data = 8'hdc;
      17'd35712: data = 8'h00;
      17'd35713: data = 8'h0e;
      17'd35714: data = 8'he9;
      17'd35715: data = 8'h06;
      17'd35716: data = 8'h05;
      17'd35717: data = 8'he9;
      17'd35718: data = 8'h00;
      17'd35719: data = 8'hfc;
      17'd35720: data = 8'hf2;
      17'd35721: data = 8'hfd;
      17'd35722: data = 8'hfe;
      17'd35723: data = 8'h0c;
      17'd35724: data = 8'hfe;
      17'd35725: data = 8'he3;
      17'd35726: data = 8'hfd;
      17'd35727: data = 8'h12;
      17'd35728: data = 8'h05;
      17'd35729: data = 8'hfd;
      17'd35730: data = 8'hf9;
      17'd35731: data = 8'hf1;
      17'd35732: data = 8'h1b;
      17'd35733: data = 8'h0e;
      17'd35734: data = 8'he7;
      17'd35735: data = 8'h02;
      17'd35736: data = 8'h09;
      17'd35737: data = 8'h06;
      17'd35738: data = 8'h16;
      17'd35739: data = 8'hf5;
      17'd35740: data = 8'hec;
      17'd35741: data = 8'h15;
      17'd35742: data = 8'h01;
      17'd35743: data = 8'h05;
      17'd35744: data = 8'hfd;
      17'd35745: data = 8'hef;
      17'd35746: data = 8'h19;
      17'd35747: data = 8'hfd;
      17'd35748: data = 8'hef;
      17'd35749: data = 8'h0a;
      17'd35750: data = 8'hfd;
      17'd35751: data = 8'h01;
      17'd35752: data = 8'hec;
      17'd35753: data = 8'h09;
      17'd35754: data = 8'h19;
      17'd35755: data = 8'he4;
      17'd35756: data = 8'hf1;
      17'd35757: data = 8'h13;
      17'd35758: data = 8'h0a;
      17'd35759: data = 8'hf1;
      17'd35760: data = 8'h00;
      17'd35761: data = 8'h0c;
      17'd35762: data = 8'h0a;
      17'd35763: data = 8'h12;
      17'd35764: data = 8'hf4;
      17'd35765: data = 8'hf2;
      17'd35766: data = 8'h24;
      17'd35767: data = 8'h0d;
      17'd35768: data = 8'hec;
      17'd35769: data = 8'h11;
      17'd35770: data = 8'h09;
      17'd35771: data = 8'hf4;
      17'd35772: data = 8'h0a;
      17'd35773: data = 8'hfe;
      17'd35774: data = 8'hf9;
      17'd35775: data = 8'h1a;
      17'd35776: data = 8'hf2;
      17'd35777: data = 8'heb;
      17'd35778: data = 8'h1e;
      17'd35779: data = 8'hf5;
      17'd35780: data = 8'he9;
      17'd35781: data = 8'h15;
      17'd35782: data = 8'h06;
      17'd35783: data = 8'hf4;
      17'd35784: data = 8'hfe;
      17'd35785: data = 8'hfe;
      17'd35786: data = 8'hfe;
      17'd35787: data = 8'h0a;
      17'd35788: data = 8'hf9;
      17'd35789: data = 8'hfe;
      17'd35790: data = 8'h0d;
      17'd35791: data = 8'hfd;
      17'd35792: data = 8'h02;
      17'd35793: data = 8'h0c;
      17'd35794: data = 8'hfa;
      17'd35795: data = 8'h04;
      17'd35796: data = 8'h01;
      17'd35797: data = 8'h04;
      17'd35798: data = 8'h0a;
      17'd35799: data = 8'hf4;
      17'd35800: data = 8'h04;
      17'd35801: data = 8'h02;
      17'd35802: data = 8'hfa;
      17'd35803: data = 8'h05;
      17'd35804: data = 8'h0c;
      17'd35805: data = 8'hf2;
      17'd35806: data = 8'hf9;
      17'd35807: data = 8'h0c;
      17'd35808: data = 8'h00;
      17'd35809: data = 8'hfe;
      17'd35810: data = 8'h01;
      17'd35811: data = 8'hf6;
      17'd35812: data = 8'heb;
      17'd35813: data = 8'h22;
      17'd35814: data = 8'h0e;
      17'd35815: data = 8'hd8;
      17'd35816: data = 8'h06;
      17'd35817: data = 8'h02;
      17'd35818: data = 8'hf4;
      17'd35819: data = 8'h1a;
      17'd35820: data = 8'h0c;
      17'd35821: data = 8'hd5;
      17'd35822: data = 8'h06;
      17'd35823: data = 8'h1a;
      17'd35824: data = 8'h00;
      17'd35825: data = 8'h04;
      17'd35826: data = 8'hed;
      17'd35827: data = 8'hfc;
      17'd35828: data = 8'h13;
      17'd35829: data = 8'h11;
      17'd35830: data = 8'hfe;
      17'd35831: data = 8'he5;
      17'd35832: data = 8'hf5;
      17'd35833: data = 8'h23;
      17'd35834: data = 8'h11;
      17'd35835: data = 8'he3;
      17'd35836: data = 8'h00;
      17'd35837: data = 8'h11;
      17'd35838: data = 8'hef;
      17'd35839: data = 8'h0d;
      17'd35840: data = 8'h09;
      17'd35841: data = 8'he4;
      17'd35842: data = 8'h1a;
      17'd35843: data = 8'h04;
      17'd35844: data = 8'heb;
      17'd35845: data = 8'h00;
      17'd35846: data = 8'hf9;
      17'd35847: data = 8'h06;
      17'd35848: data = 8'hf4;
      17'd35849: data = 8'hf4;
      17'd35850: data = 8'h0a;
      17'd35851: data = 8'he5;
      17'd35852: data = 8'hf5;
      17'd35853: data = 8'h12;
      17'd35854: data = 8'he7;
      17'd35855: data = 8'hfc;
      17'd35856: data = 8'h0e;
      17'd35857: data = 8'he3;
      17'd35858: data = 8'h11;
      17'd35859: data = 8'h0e;
      17'd35860: data = 8'hd8;
      17'd35861: data = 8'h09;
      17'd35862: data = 8'h23;
      17'd35863: data = 8'hf5;
      17'd35864: data = 8'hf4;
      17'd35865: data = 8'h04;
      17'd35866: data = 8'hf5;
      17'd35867: data = 8'h06;
      17'd35868: data = 8'h1a;
      17'd35869: data = 8'h02;
      17'd35870: data = 8'hed;
      17'd35871: data = 8'hf2;
      17'd35872: data = 8'h0a;
      17'd35873: data = 8'h05;
      17'd35874: data = 8'h01;
      17'd35875: data = 8'hfd;
      17'd35876: data = 8'hed;
      17'd35877: data = 8'h01;
      17'd35878: data = 8'hfd;
      17'd35879: data = 8'h05;
      17'd35880: data = 8'h02;
      17'd35881: data = 8'hec;
      17'd35882: data = 8'hfe;
      17'd35883: data = 8'h00;
      17'd35884: data = 8'h0a;
      17'd35885: data = 8'hfa;
      17'd35886: data = 8'he7;
      17'd35887: data = 8'h12;
      17'd35888: data = 8'h04;
      17'd35889: data = 8'heb;
      17'd35890: data = 8'h04;
      17'd35891: data = 8'h00;
      17'd35892: data = 8'hf1;
      17'd35893: data = 8'h0e;
      17'd35894: data = 8'h02;
      17'd35895: data = 8'hef;
      17'd35896: data = 8'h00;
      17'd35897: data = 8'h0a;
      17'd35898: data = 8'h04;
      17'd35899: data = 8'hf6;
      17'd35900: data = 8'h0a;
      17'd35901: data = 8'h00;
      17'd35902: data = 8'he2;
      17'd35903: data = 8'h24;
      17'd35904: data = 8'h09;
      17'd35905: data = 8'hd8;
      17'd35906: data = 8'h0c;
      17'd35907: data = 8'h05;
      17'd35908: data = 8'hfa;
      17'd35909: data = 8'hfd;
      17'd35910: data = 8'hf9;
      17'd35911: data = 8'hfc;
      17'd35912: data = 8'hfa;
      17'd35913: data = 8'h09;
      17'd35914: data = 8'h00;
      17'd35915: data = 8'he7;
      17'd35916: data = 8'h11;
      17'd35917: data = 8'h11;
      17'd35918: data = 8'hec;
      17'd35919: data = 8'hfd;
      17'd35920: data = 8'h0e;
      17'd35921: data = 8'hf5;
      17'd35922: data = 8'hf2;
      17'd35923: data = 8'h1b;
      17'd35924: data = 8'h02;
      17'd35925: data = 8'he5;
      17'd35926: data = 8'h04;
      17'd35927: data = 8'hfc;
      17'd35928: data = 8'hfc;
      17'd35929: data = 8'h0a;
      17'd35930: data = 8'hfa;
      17'd35931: data = 8'he4;
      17'd35932: data = 8'hfc;
      17'd35933: data = 8'h12;
      17'd35934: data = 8'h02;
      17'd35935: data = 8'hed;
      17'd35936: data = 8'hf9;
      17'd35937: data = 8'h0d;
      17'd35938: data = 8'hf6;
      17'd35939: data = 8'h0e;
      17'd35940: data = 8'h06;
      17'd35941: data = 8'he7;
      17'd35942: data = 8'h09;
      17'd35943: data = 8'h06;
      17'd35944: data = 8'hf9;
      17'd35945: data = 8'h11;
      17'd35946: data = 8'h04;
      17'd35947: data = 8'hec;
      17'd35948: data = 8'hf4;
      17'd35949: data = 8'h04;
      17'd35950: data = 8'h13;
      17'd35951: data = 8'hef;
      17'd35952: data = 8'he9;
      17'd35953: data = 8'h22;
      17'd35954: data = 8'he0;
      17'd35955: data = 8'hdc;
      17'd35956: data = 8'h2c;
      17'd35957: data = 8'hfa;
      17'd35958: data = 8'hed;
      17'd35959: data = 8'h06;
      17'd35960: data = 8'he0;
      17'd35961: data = 8'h01;
      17'd35962: data = 8'h2f;
      17'd35963: data = 8'he9;
      17'd35964: data = 8'he0;
      17'd35965: data = 8'h15;
      17'd35966: data = 8'h0d;
      17'd35967: data = 8'h05;
      17'd35968: data = 8'h05;
      17'd35969: data = 8'hf6;
      17'd35970: data = 8'he9;
      17'd35971: data = 8'h12;
      17'd35972: data = 8'h33;
      17'd35973: data = 8'hf9;
      17'd35974: data = 8'hde;
      17'd35975: data = 8'hf4;
      17'd35976: data = 8'h0c;
      17'd35977: data = 8'h15;
      17'd35978: data = 8'h1b;
      17'd35979: data = 8'hec;
      17'd35980: data = 8'hd8;
      17'd35981: data = 8'h0e;
      17'd35982: data = 8'h27;
      17'd35983: data = 8'h12;
      17'd35984: data = 8'hdb;
      17'd35985: data = 8'hfa;
      17'd35986: data = 8'h09;
      17'd35987: data = 8'h0a;
      17'd35988: data = 8'h11;
      17'd35989: data = 8'he3;
      17'd35990: data = 8'hfa;
      17'd35991: data = 8'hf9;
      17'd35992: data = 8'h1e;
      17'd35993: data = 8'h1b;
      17'd35994: data = 8'hc4;
      17'd35995: data = 8'hfa;
      17'd35996: data = 8'h22;
      17'd35997: data = 8'hfc;
      17'd35998: data = 8'h1b;
      17'd35999: data = 8'hef;
      17'd36000: data = 8'hd2;
      17'd36001: data = 8'h1c;
      17'd36002: data = 8'h24;
      17'd36003: data = 8'h06;
      17'd36004: data = 8'hf2;
      17'd36005: data = 8'hec;
      17'd36006: data = 8'hf2;
      17'd36007: data = 8'h24;
      17'd36008: data = 8'h1a;
      17'd36009: data = 8'hed;
      17'd36010: data = 8'hfd;
      17'd36011: data = 8'heb;
      17'd36012: data = 8'h0e;
      17'd36013: data = 8'h35;
      17'd36014: data = 8'he3;
      17'd36015: data = 8'hd8;
      17'd36016: data = 8'h19;
      17'd36017: data = 8'h12;
      17'd36018: data = 8'h09;
      17'd36019: data = 8'hf6;
      17'd36020: data = 8'he3;
      17'd36021: data = 8'hfa;
      17'd36022: data = 8'h1e;
      17'd36023: data = 8'h16;
      17'd36024: data = 8'he3;
      17'd36025: data = 8'hed;
      17'd36026: data = 8'h13;
      17'd36027: data = 8'hfc;
      17'd36028: data = 8'h02;
      17'd36029: data = 8'h1b;
      17'd36030: data = 8'he2;
      17'd36031: data = 8'hec;
      17'd36032: data = 8'h22;
      17'd36033: data = 8'h0a;
      17'd36034: data = 8'hed;
      17'd36035: data = 8'hf2;
      17'd36036: data = 8'h00;
      17'd36037: data = 8'h05;
      17'd36038: data = 8'h0c;
      17'd36039: data = 8'h01;
      17'd36040: data = 8'hed;
      17'd36041: data = 8'hf6;
      17'd36042: data = 8'h19;
      17'd36043: data = 8'h09;
      17'd36044: data = 8'hf1;
      17'd36045: data = 8'h1c;
      17'd36046: data = 8'h0c;
      17'd36047: data = 8'hd8;
      17'd36048: data = 8'h0a;
      17'd36049: data = 8'h19;
      17'd36050: data = 8'hfc;
      17'd36051: data = 8'hf6;
      17'd36052: data = 8'h0a;
      17'd36053: data = 8'hf5;
      17'd36054: data = 8'he9;
      17'd36055: data = 8'h05;
      17'd36056: data = 8'h0a;
      17'd36057: data = 8'h02;
      17'd36058: data = 8'hf1;
      17'd36059: data = 8'hf1;
      17'd36060: data = 8'hfd;
      17'd36061: data = 8'h04;
      17'd36062: data = 8'h06;
      17'd36063: data = 8'hfa;
      17'd36064: data = 8'hfa;
      17'd36065: data = 8'hfe;
      17'd36066: data = 8'h02;
      17'd36067: data = 8'h01;
      17'd36068: data = 8'hfc;
      17'd36069: data = 8'h0e;
      17'd36070: data = 8'h02;
      17'd36071: data = 8'hec;
      17'd36072: data = 8'hfc;
      17'd36073: data = 8'h12;
      17'd36074: data = 8'h1a;
      17'd36075: data = 8'hf5;
      17'd36076: data = 8'he5;
      17'd36077: data = 8'h0a;
      17'd36078: data = 8'h15;
      17'd36079: data = 8'h09;
      17'd36080: data = 8'hf6;
      17'd36081: data = 8'hfa;
      17'd36082: data = 8'hfa;
      17'd36083: data = 8'h00;
      17'd36084: data = 8'h13;
      17'd36085: data = 8'hf1;
      17'd36086: data = 8'hf4;
      17'd36087: data = 8'h01;
      17'd36088: data = 8'heb;
      17'd36089: data = 8'hfe;
      17'd36090: data = 8'h13;
      17'd36091: data = 8'hdb;
      17'd36092: data = 8'hf1;
      17'd36093: data = 8'h1b;
      17'd36094: data = 8'hda;
      17'd36095: data = 8'h02;
      17'd36096: data = 8'h0c;
      17'd36097: data = 8'he2;
      17'd36098: data = 8'h0e;
      17'd36099: data = 8'hfd;
      17'd36100: data = 8'h04;
      17'd36101: data = 8'h0d;
      17'd36102: data = 8'hef;
      17'd36103: data = 8'h1f;
      17'd36104: data = 8'h01;
      17'd36105: data = 8'hed;
      17'd36106: data = 8'h0c;
      17'd36107: data = 8'h2b;
      17'd36108: data = 8'h11;
      17'd36109: data = 8'hcb;
      17'd36110: data = 8'h09;
      17'd36111: data = 8'h12;
      17'd36112: data = 8'hef;
      17'd36113: data = 8'h1a;
      17'd36114: data = 8'hf6;
      17'd36115: data = 8'he0;
      17'd36116: data = 8'h04;
      17'd36117: data = 8'h04;
      17'd36118: data = 8'hfd;
      17'd36119: data = 8'hf9;
      17'd36120: data = 8'hf9;
      17'd36121: data = 8'hfa;
      17'd36122: data = 8'h0c;
      17'd36123: data = 8'hf1;
      17'd36124: data = 8'heb;
      17'd36125: data = 8'h12;
      17'd36126: data = 8'h04;
      17'd36127: data = 8'hf2;
      17'd36128: data = 8'h0a;
      17'd36129: data = 8'hf4;
      17'd36130: data = 8'hfa;
      17'd36131: data = 8'h19;
      17'd36132: data = 8'heb;
      17'd36133: data = 8'heb;
      17'd36134: data = 8'h1a;
      17'd36135: data = 8'h12;
      17'd36136: data = 8'hef;
      17'd36137: data = 8'h11;
      17'd36138: data = 8'heb;
      17'd36139: data = 8'he7;
      17'd36140: data = 8'h34;
      17'd36141: data = 8'hf9;
      17'd36142: data = 8'he4;
      17'd36143: data = 8'h1b;
      17'd36144: data = 8'he7;
      17'd36145: data = 8'hf5;
      17'd36146: data = 8'h1c;
      17'd36147: data = 8'hed;
      17'd36148: data = 8'hf6;
      17'd36149: data = 8'h09;
      17'd36150: data = 8'hf5;
      17'd36151: data = 8'h01;
      17'd36152: data = 8'h15;
      17'd36153: data = 8'hd8;
      17'd36154: data = 8'hfa;
      17'd36155: data = 8'h29;
      17'd36156: data = 8'he9;
      17'd36157: data = 8'hfa;
      17'd36158: data = 8'h04;
      17'd36159: data = 8'hec;
      17'd36160: data = 8'h05;
      17'd36161: data = 8'h1f;
      17'd36162: data = 8'he7;
      17'd36163: data = 8'he4;
      17'd36164: data = 8'h24;
      17'd36165: data = 8'hf5;
      17'd36166: data = 8'hf2;
      17'd36167: data = 8'h11;
      17'd36168: data = 8'hf4;
      17'd36169: data = 8'hf4;
      17'd36170: data = 8'h02;
      17'd36171: data = 8'hf9;
      17'd36172: data = 8'h05;
      17'd36173: data = 8'h05;
      17'd36174: data = 8'hf6;
      17'd36175: data = 8'h09;
      17'd36176: data = 8'hf9;
      17'd36177: data = 8'hf6;
      17'd36178: data = 8'h0e;
      17'd36179: data = 8'hfa;
      17'd36180: data = 8'h01;
      17'd36181: data = 8'h1b;
      17'd36182: data = 8'he7;
      17'd36183: data = 8'he5;
      17'd36184: data = 8'h15;
      17'd36185: data = 8'h0e;
      17'd36186: data = 8'hf9;
      17'd36187: data = 8'hef;
      17'd36188: data = 8'he2;
      17'd36189: data = 8'h04;
      17'd36190: data = 8'h2c;
      17'd36191: data = 8'he3;
      17'd36192: data = 8'hd2;
      17'd36193: data = 8'h16;
      17'd36194: data = 8'h02;
      17'd36195: data = 8'hf6;
      17'd36196: data = 8'h05;
      17'd36197: data = 8'he5;
      17'd36198: data = 8'hf9;
      17'd36199: data = 8'h12;
      17'd36200: data = 8'h04;
      17'd36201: data = 8'h05;
      17'd36202: data = 8'hf2;
      17'd36203: data = 8'hf5;
      17'd36204: data = 8'h05;
      17'd36205: data = 8'h22;
      17'd36206: data = 8'h13;
      17'd36207: data = 8'hd5;
      17'd36208: data = 8'h00;
      17'd36209: data = 8'h12;
      17'd36210: data = 8'h12;
      17'd36211: data = 8'h12;
      17'd36212: data = 8'hcb;
      17'd36213: data = 8'hf9;
      17'd36214: data = 8'h27;
      17'd36215: data = 8'hf6;
      17'd36216: data = 8'h02;
      17'd36217: data = 8'h00;
      17'd36218: data = 8'he2;
      17'd36219: data = 8'h0d;
      17'd36220: data = 8'h1f;
      17'd36221: data = 8'hef;
      17'd36222: data = 8'he7;
      17'd36223: data = 8'h00;
      17'd36224: data = 8'h09;
      17'd36225: data = 8'h05;
      17'd36226: data = 8'hfe;
      17'd36227: data = 8'heb;
      17'd36228: data = 8'he7;
      17'd36229: data = 8'h1f;
      17'd36230: data = 8'h0d;
      17'd36231: data = 8'hde;
      17'd36232: data = 8'hf1;
      17'd36233: data = 8'h05;
      17'd36234: data = 8'h1a;
      17'd36235: data = 8'hfd;
      17'd36236: data = 8'h01;
      17'd36237: data = 8'hfc;
      17'd36238: data = 8'hde;
      17'd36239: data = 8'h1c;
      17'd36240: data = 8'h1e;
      17'd36241: data = 8'he9;
      17'd36242: data = 8'hfa;
      17'd36243: data = 8'h01;
      17'd36244: data = 8'h01;
      17'd36245: data = 8'h0e;
      17'd36246: data = 8'h0c;
      17'd36247: data = 8'he5;
      17'd36248: data = 8'hec;
      17'd36249: data = 8'h1e;
      17'd36250: data = 8'h05;
      17'd36251: data = 8'hef;
      17'd36252: data = 8'h06;
      17'd36253: data = 8'hfc;
      17'd36254: data = 8'hf5;
      17'd36255: data = 8'h09;
      17'd36256: data = 8'hf9;
      17'd36257: data = 8'h0e;
      17'd36258: data = 8'hef;
      17'd36259: data = 8'he4;
      17'd36260: data = 8'h19;
      17'd36261: data = 8'h04;
      17'd36262: data = 8'hf4;
      17'd36263: data = 8'hef;
      17'd36264: data = 8'h15;
      17'd36265: data = 8'hf1;
      17'd36266: data = 8'hfc;
      17'd36267: data = 8'h2c;
      17'd36268: data = 8'hd5;
      17'd36269: data = 8'hf2;
      17'd36270: data = 8'h2f;
      17'd36271: data = 8'hf4;
      17'd36272: data = 8'hf5;
      17'd36273: data = 8'h0a;
      17'd36274: data = 8'hf4;
      17'd36275: data = 8'h0a;
      17'd36276: data = 8'h15;
      17'd36277: data = 8'hed;
      17'd36278: data = 8'h04;
      17'd36279: data = 8'h00;
      17'd36280: data = 8'hf1;
      17'd36281: data = 8'h23;
      17'd36282: data = 8'h0a;
      17'd36283: data = 8'hd8;
      17'd36284: data = 8'hfc;
      17'd36285: data = 8'h0c;
      17'd36286: data = 8'hf9;
      17'd36287: data = 8'h0c;
      17'd36288: data = 8'hfc;
      17'd36289: data = 8'he3;
      17'd36290: data = 8'hfe;
      17'd36291: data = 8'hfe;
      17'd36292: data = 8'hfe;
      17'd36293: data = 8'hfa;
      17'd36294: data = 8'hf6;
      17'd36295: data = 8'h04;
      17'd36296: data = 8'hec;
      17'd36297: data = 8'h01;
      17'd36298: data = 8'hfe;
      17'd36299: data = 8'hf4;
      17'd36300: data = 8'h06;
      17'd36301: data = 8'hf2;
      17'd36302: data = 8'h15;
      17'd36303: data = 8'h05;
      17'd36304: data = 8'he9;
      17'd36305: data = 8'h15;
      17'd36306: data = 8'hfd;
      17'd36307: data = 8'h09;
      17'd36308: data = 8'h19;
      17'd36309: data = 8'hf2;
      17'd36310: data = 8'h02;
      17'd36311: data = 8'h13;
      17'd36312: data = 8'h00;
      17'd36313: data = 8'hf2;
      17'd36314: data = 8'h02;
      17'd36315: data = 8'h02;
      17'd36316: data = 8'hfd;
      17'd36317: data = 8'h16;
      17'd36318: data = 8'hec;
      17'd36319: data = 8'he7;
      17'd36320: data = 8'h1b;
      17'd36321: data = 8'hf2;
      17'd36322: data = 8'hf2;
      17'd36323: data = 8'h09;
      17'd36324: data = 8'hed;
      17'd36325: data = 8'h01;
      17'd36326: data = 8'hf6;
      17'd36327: data = 8'hdc;
      17'd36328: data = 8'h1b;
      17'd36329: data = 8'hfd;
      17'd36330: data = 8'hdc;
      17'd36331: data = 8'h11;
      17'd36332: data = 8'hfd;
      17'd36333: data = 8'hfa;
      17'd36334: data = 8'h05;
      17'd36335: data = 8'hf5;
      17'd36336: data = 8'h11;
      17'd36337: data = 8'h01;
      17'd36338: data = 8'hfa;
      17'd36339: data = 8'h12;
      17'd36340: data = 8'hfd;
      17'd36341: data = 8'h0c;
      17'd36342: data = 8'h00;
      17'd36343: data = 8'hf9;
      17'd36344: data = 8'h02;
      17'd36345: data = 8'h0d;
      17'd36346: data = 8'h0a;
      17'd36347: data = 8'hde;
      17'd36348: data = 8'h13;
      17'd36349: data = 8'h11;
      17'd36350: data = 8'hde;
      17'd36351: data = 8'h0e;
      17'd36352: data = 8'hfa;
      17'd36353: data = 8'hf1;
      17'd36354: data = 8'h16;
      17'd36355: data = 8'hed;
      17'd36356: data = 8'hf5;
      17'd36357: data = 8'h02;
      17'd36358: data = 8'hed;
      17'd36359: data = 8'h05;
      17'd36360: data = 8'h04;
      17'd36361: data = 8'hf9;
      17'd36362: data = 8'hfc;
      17'd36363: data = 8'hf5;
      17'd36364: data = 8'h0c;
      17'd36365: data = 8'hfa;
      17'd36366: data = 8'hfe;
      17'd36367: data = 8'h0d;
      17'd36368: data = 8'hec;
      17'd36369: data = 8'h16;
      17'd36370: data = 8'hfd;
      17'd36371: data = 8'hed;
      17'd36372: data = 8'h23;
      17'd36373: data = 8'hf6;
      17'd36374: data = 8'hf5;
      17'd36375: data = 8'h11;
      17'd36376: data = 8'hfc;
      17'd36377: data = 8'h05;
      17'd36378: data = 8'h00;
      17'd36379: data = 8'hf6;
      17'd36380: data = 8'h04;
      17'd36381: data = 8'hed;
      17'd36382: data = 8'h01;
      17'd36383: data = 8'h0c;
      17'd36384: data = 8'he9;
      17'd36385: data = 8'hfe;
      17'd36386: data = 8'h06;
      17'd36387: data = 8'hf2;
      17'd36388: data = 8'hf9;
      17'd36389: data = 8'h04;
      17'd36390: data = 8'h00;
      17'd36391: data = 8'h04;
      17'd36392: data = 8'hfd;
      17'd36393: data = 8'hf1;
      17'd36394: data = 8'h05;
      17'd36395: data = 8'h0c;
      17'd36396: data = 8'hfe;
      17'd36397: data = 8'hfe;
      17'd36398: data = 8'h04;
      17'd36399: data = 8'hed;
      17'd36400: data = 8'hfd;
      17'd36401: data = 8'h09;
      17'd36402: data = 8'hfc;
      17'd36403: data = 8'h00;
      17'd36404: data = 8'hf4;
      17'd36405: data = 8'hfe;
      17'd36406: data = 8'h00;
      17'd36407: data = 8'h04;
      17'd36408: data = 8'h02;
      17'd36409: data = 8'heb;
      17'd36410: data = 8'h02;
      17'd36411: data = 8'h1b;
      17'd36412: data = 8'hf9;
      17'd36413: data = 8'hf6;
      17'd36414: data = 8'h09;
      17'd36415: data = 8'hf9;
      17'd36416: data = 8'hfe;
      17'd36417: data = 8'h04;
      17'd36418: data = 8'hfd;
      17'd36419: data = 8'h05;
      17'd36420: data = 8'hf5;
      17'd36421: data = 8'hf4;
      17'd36422: data = 8'h04;
      17'd36423: data = 8'hfe;
      17'd36424: data = 8'h02;
      17'd36425: data = 8'hf2;
      17'd36426: data = 8'hf5;
      17'd36427: data = 8'h09;
      17'd36428: data = 8'hfa;
      17'd36429: data = 8'hf9;
      17'd36430: data = 8'h06;
      17'd36431: data = 8'h04;
      17'd36432: data = 8'hf4;
      17'd36433: data = 8'h0a;
      17'd36434: data = 8'h0c;
      17'd36435: data = 8'hec;
      17'd36436: data = 8'h04;
      17'd36437: data = 8'h12;
      17'd36438: data = 8'hfe;
      17'd36439: data = 8'h05;
      17'd36440: data = 8'h02;
      17'd36441: data = 8'hfe;
      17'd36442: data = 8'h0c;
      17'd36443: data = 8'hfc;
      17'd36444: data = 8'hfc;
      17'd36445: data = 8'h04;
      17'd36446: data = 8'hfa;
      17'd36447: data = 8'h00;
      17'd36448: data = 8'h0c;
      17'd36449: data = 8'hfc;
      17'd36450: data = 8'hf5;
      17'd36451: data = 8'h01;
      17'd36452: data = 8'h00;
      17'd36453: data = 8'h02;
      17'd36454: data = 8'h0a;
      17'd36455: data = 8'h00;
      17'd36456: data = 8'hf5;
      17'd36457: data = 8'h00;
      17'd36458: data = 8'h05;
      17'd36459: data = 8'h00;
      17'd36460: data = 8'hfe;
      17'd36461: data = 8'hfc;
      17'd36462: data = 8'h02;
      17'd36463: data = 8'hfe;
      17'd36464: data = 8'hf9;
      17'd36465: data = 8'h04;
      17'd36466: data = 8'h02;
      17'd36467: data = 8'hfa;
      17'd36468: data = 8'h05;
      17'd36469: data = 8'h01;
      17'd36470: data = 8'h01;
      17'd36471: data = 8'h0c;
      17'd36472: data = 8'hfd;
      17'd36473: data = 8'hf6;
      17'd36474: data = 8'h05;
      17'd36475: data = 8'h0d;
      17'd36476: data = 8'hfc;
      17'd36477: data = 8'h00;
      17'd36478: data = 8'h09;
      17'd36479: data = 8'hf4;
      17'd36480: data = 8'hfd;
      17'd36481: data = 8'h0e;
      17'd36482: data = 8'h05;
      17'd36483: data = 8'h01;
      17'd36484: data = 8'hf9;
      17'd36485: data = 8'hfd;
      17'd36486: data = 8'h05;
      17'd36487: data = 8'h06;
      17'd36488: data = 8'h02;
      17'd36489: data = 8'hef;
      17'd36490: data = 8'hfc;
      17'd36491: data = 8'h0c;
      17'd36492: data = 8'hfe;
      17'd36493: data = 8'hfa;
      17'd36494: data = 8'h00;
      17'd36495: data = 8'hfc;
      17'd36496: data = 8'h04;
      17'd36497: data = 8'h04;
      17'd36498: data = 8'hf4;
      17'd36499: data = 8'h04;
      17'd36500: data = 8'h02;
      17'd36501: data = 8'hf5;
      17'd36502: data = 8'h02;
      17'd36503: data = 8'h01;
      17'd36504: data = 8'hf2;
      17'd36505: data = 8'hfa;
      17'd36506: data = 8'hfa;
      17'd36507: data = 8'hfc;
      17'd36508: data = 8'h0c;
      17'd36509: data = 8'hf5;
      17'd36510: data = 8'hf1;
      17'd36511: data = 8'h0a;
      17'd36512: data = 8'h02;
      17'd36513: data = 8'hfa;
      17'd36514: data = 8'h01;
      17'd36515: data = 8'h00;
      17'd36516: data = 8'h05;
      17'd36517: data = 8'h01;
      17'd36518: data = 8'hf2;
      17'd36519: data = 8'h02;
      17'd36520: data = 8'h02;
      17'd36521: data = 8'hfd;
      17'd36522: data = 8'hfa;
      17'd36523: data = 8'hf1;
      17'd36524: data = 8'h09;
      17'd36525: data = 8'h05;
      17'd36526: data = 8'hf2;
      17'd36527: data = 8'h01;
      17'd36528: data = 8'hfd;
      17'd36529: data = 8'hf9;
      17'd36530: data = 8'h02;
      17'd36531: data = 8'hf9;
      17'd36532: data = 8'hf9;
      17'd36533: data = 8'h04;
      17'd36534: data = 8'hfe;
      17'd36535: data = 8'hf6;
      17'd36536: data = 8'hfc;
      17'd36537: data = 8'h01;
      17'd36538: data = 8'h01;
      17'd36539: data = 8'h00;
      17'd36540: data = 8'h02;
      17'd36541: data = 8'h05;
      17'd36542: data = 8'hfd;
      17'd36543: data = 8'hfd;
      17'd36544: data = 8'h00;
      17'd36545: data = 8'h06;
      17'd36546: data = 8'h02;
      17'd36547: data = 8'hfc;
      17'd36548: data = 8'hfe;
      17'd36549: data = 8'hfc;
      17'd36550: data = 8'h02;
      17'd36551: data = 8'h01;
      17'd36552: data = 8'hf2;
      17'd36553: data = 8'h04;
      17'd36554: data = 8'h09;
      17'd36555: data = 8'h02;
      17'd36556: data = 8'hfc;
      17'd36557: data = 8'hed;
      17'd36558: data = 8'h05;
      17'd36559: data = 8'h06;
      17'd36560: data = 8'hfe;
      17'd36561: data = 8'h00;
      17'd36562: data = 8'heb;
      17'd36563: data = 8'hfc;
      17'd36564: data = 8'h04;
      17'd36565: data = 8'hf2;
      17'd36566: data = 8'h01;
      17'd36567: data = 8'h01;
      17'd36568: data = 8'hf4;
      17'd36569: data = 8'hf9;
      17'd36570: data = 8'hfe;
      17'd36571: data = 8'h09;
      17'd36572: data = 8'h05;
      17'd36573: data = 8'h01;
      17'd36574: data = 8'h04;
      17'd36575: data = 8'hfd;
      17'd36576: data = 8'h04;
      17'd36577: data = 8'h09;
      17'd36578: data = 8'h02;
      17'd36579: data = 8'h0a;
      17'd36580: data = 8'h00;
      17'd36581: data = 8'hf5;
      17'd36582: data = 8'h00;
      17'd36583: data = 8'h0d;
      17'd36584: data = 8'h00;
      17'd36585: data = 8'hf4;
      17'd36586: data = 8'h01;
      17'd36587: data = 8'hf6;
      17'd36588: data = 8'hfe;
      17'd36589: data = 8'h06;
      17'd36590: data = 8'hf5;
      17'd36591: data = 8'h04;
      17'd36592: data = 8'h00;
      17'd36593: data = 8'hfd;
      17'd36594: data = 8'h06;
      17'd36595: data = 8'hfa;
      17'd36596: data = 8'h02;
      17'd36597: data = 8'hfd;
      17'd36598: data = 8'h00;
      17'd36599: data = 8'h13;
      17'd36600: data = 8'hf9;
      17'd36601: data = 8'hf5;
      17'd36602: data = 8'h02;
      17'd36603: data = 8'hfd;
      17'd36604: data = 8'h05;
      17'd36605: data = 8'h09;
      17'd36606: data = 8'hfd;
      17'd36607: data = 8'hf5;
      17'd36608: data = 8'hfe;
      17'd36609: data = 8'h0a;
      17'd36610: data = 8'h02;
      17'd36611: data = 8'h0a;
      17'd36612: data = 8'h00;
      17'd36613: data = 8'hf2;
      17'd36614: data = 8'h0a;
      17'd36615: data = 8'h04;
      17'd36616: data = 8'h06;
      17'd36617: data = 8'h00;
      17'd36618: data = 8'hf4;
      17'd36619: data = 8'h0c;
      17'd36620: data = 8'h0a;
      17'd36621: data = 8'hf1;
      17'd36622: data = 8'hfa;
      17'd36623: data = 8'h09;
      17'd36624: data = 8'hf6;
      17'd36625: data = 8'hfd;
      17'd36626: data = 8'hfd;
      17'd36627: data = 8'hf4;
      17'd36628: data = 8'h04;
      17'd36629: data = 8'h01;
      17'd36630: data = 8'hfd;
      17'd36631: data = 8'h00;
      17'd36632: data = 8'hfe;
      17'd36633: data = 8'hfe;
      17'd36634: data = 8'h06;
      17'd36635: data = 8'h05;
      17'd36636: data = 8'hf9;
      17'd36637: data = 8'hfe;
      17'd36638: data = 8'h01;
      17'd36639: data = 8'h04;
      17'd36640: data = 8'h05;
      17'd36641: data = 8'hf9;
      17'd36642: data = 8'hf5;
      17'd36643: data = 8'h00;
      17'd36644: data = 8'h06;
      17'd36645: data = 8'h02;
      17'd36646: data = 8'hfc;
      17'd36647: data = 8'hfd;
      17'd36648: data = 8'h01;
      17'd36649: data = 8'h06;
      17'd36650: data = 8'h05;
      17'd36651: data = 8'hfd;
      17'd36652: data = 8'hfe;
      17'd36653: data = 8'h00;
      17'd36654: data = 8'hfd;
      17'd36655: data = 8'h05;
      17'd36656: data = 8'h01;
      17'd36657: data = 8'hfa;
      17'd36658: data = 8'h00;
      17'd36659: data = 8'hfe;
      17'd36660: data = 8'hfd;
      17'd36661: data = 8'h00;
      17'd36662: data = 8'h00;
      17'd36663: data = 8'h00;
      17'd36664: data = 8'h00;
      17'd36665: data = 8'h00;
      17'd36666: data = 8'h00;
      17'd36667: data = 8'h02;
      17'd36668: data = 8'h01;
      17'd36669: data = 8'h01;
      17'd36670: data = 8'h01;
      17'd36671: data = 8'hfe;
      17'd36672: data = 8'h00;
      17'd36673: data = 8'h01;
      17'd36674: data = 8'h01;
      17'd36675: data = 8'h01;
      17'd36676: data = 8'h01;
      17'd36677: data = 8'h01;
      17'd36678: data = 8'h00;
      17'd36679: data = 8'hfe;
      17'd36680: data = 8'h01;
      17'd36681: data = 8'h00;
      17'd36682: data = 8'hfc;
      17'd36683: data = 8'h00;
      17'd36684: data = 8'h01;
      17'd36685: data = 8'hfe;
      17'd36686: data = 8'h01;
      17'd36687: data = 8'h04;
      17'd36688: data = 8'h02;
      17'd36689: data = 8'h04;
      17'd36690: data = 8'h02;
      17'd36691: data = 8'hfe;
      17'd36692: data = 8'h02;
      17'd36693: data = 8'h04;
      17'd36694: data = 8'h05;
      17'd36695: data = 8'h02;
      17'd36696: data = 8'hfe;
      17'd36697: data = 8'hfd;
      17'd36698: data = 8'hfd;
      17'd36699: data = 8'h01;
      17'd36700: data = 8'h01;
      17'd36701: data = 8'hfc;
      17'd36702: data = 8'hfa;
      17'd36703: data = 8'hfd;
      17'd36704: data = 8'h05;
      17'd36705: data = 8'h02;
      17'd36706: data = 8'h00;
      17'd36707: data = 8'h00;
      17'd36708: data = 8'h02;
      17'd36709: data = 8'h01;
      17'd36710: data = 8'h00;
      17'd36711: data = 8'h05;
      17'd36712: data = 8'h01;
      17'd36713: data = 8'h00;
      17'd36714: data = 8'h00;
      17'd36715: data = 8'hfc;
      17'd36716: data = 8'h01;
      17'd36717: data = 8'h04;
      17'd36718: data = 8'hfa;
      17'd36719: data = 8'hfa;
      17'd36720: data = 8'h01;
      17'd36721: data = 8'h00;
      17'd36722: data = 8'h04;
      17'd36723: data = 8'h02;
      17'd36724: data = 8'hfd;
      17'd36725: data = 8'h01;
      17'd36726: data = 8'hfd;
      17'd36727: data = 8'hfe;
      17'd36728: data = 8'h04;
      17'd36729: data = 8'h00;
      17'd36730: data = 8'hfa;
      17'd36731: data = 8'hf6;
      17'd36732: data = 8'hfa;
      17'd36733: data = 8'h02;
      17'd36734: data = 8'hfd;
      17'd36735: data = 8'hfd;
      17'd36736: data = 8'hfc;
      17'd36737: data = 8'hf9;
      17'd36738: data = 8'hfe;
      17'd36739: data = 8'hfd;
      17'd36740: data = 8'h00;
      17'd36741: data = 8'hfd;
      17'd36742: data = 8'h00;
      17'd36743: data = 8'h00;
      17'd36744: data = 8'hfa;
      17'd36745: data = 8'hfc;
      17'd36746: data = 8'hfd;
      17'd36747: data = 8'h04;
      17'd36748: data = 8'h02;
      17'd36749: data = 8'hfc;
      17'd36750: data = 8'h05;
      17'd36751: data = 8'h09;
      17'd36752: data = 8'hfc;
      17'd36753: data = 8'h04;
      17'd36754: data = 8'h00;
      17'd36755: data = 8'h04;
      17'd36756: data = 8'h09;
      17'd36757: data = 8'hfd;
      17'd36758: data = 8'h01;
      17'd36759: data = 8'h00;
      17'd36760: data = 8'hfd;
      17'd36761: data = 8'h01;
      17'd36762: data = 8'h01;
      17'd36763: data = 8'hfa;
      17'd36764: data = 8'hfa;
      17'd36765: data = 8'h01;
      17'd36766: data = 8'hfd;
      17'd36767: data = 8'hfe;
      17'd36768: data = 8'h00;
      17'd36769: data = 8'hfc;
      17'd36770: data = 8'h02;
      17'd36771: data = 8'hfe;
      17'd36772: data = 8'h00;
      17'd36773: data = 8'h01;
      17'd36774: data = 8'hf4;
      17'd36775: data = 8'h02;
      17'd36776: data = 8'h06;
      17'd36777: data = 8'hf9;
      17'd36778: data = 8'hfe;
      17'd36779: data = 8'h04;
      17'd36780: data = 8'hfd;
      17'd36781: data = 8'h01;
      17'd36782: data = 8'h04;
      17'd36783: data = 8'hfd;
      17'd36784: data = 8'h05;
      17'd36785: data = 8'h04;
      17'd36786: data = 8'hfd;
      17'd36787: data = 8'h01;
      17'd36788: data = 8'h00;
      17'd36789: data = 8'hfd;
      17'd36790: data = 8'h00;
      17'd36791: data = 8'h00;
      17'd36792: data = 8'hfd;
      17'd36793: data = 8'hfa;
      17'd36794: data = 8'hfd;
      17'd36795: data = 8'hfa;
      17'd36796: data = 8'h01;
      17'd36797: data = 8'hfe;
      17'd36798: data = 8'hfc;
      17'd36799: data = 8'hfd;
      17'd36800: data = 8'hf9;
      17'd36801: data = 8'hfd;
      17'd36802: data = 8'hfd;
      17'd36803: data = 8'hfa;
      17'd36804: data = 8'hfa;
      17'd36805: data = 8'hfc;
      17'd36806: data = 8'hfa;
      17'd36807: data = 8'hfc;
      17'd36808: data = 8'h00;
      17'd36809: data = 8'hfd;
      17'd36810: data = 8'hfd;
      17'd36811: data = 8'h01;
      17'd36812: data = 8'h01;
      17'd36813: data = 8'h00;
      17'd36814: data = 8'h02;
      17'd36815: data = 8'hfe;
      17'd36816: data = 8'h02;
      17'd36817: data = 8'h05;
      17'd36818: data = 8'h01;
      17'd36819: data = 8'hfe;
      17'd36820: data = 8'hfe;
      17'd36821: data = 8'hfe;
      17'd36822: data = 8'h01;
      17'd36823: data = 8'h00;
      17'd36824: data = 8'hf9;
      17'd36825: data = 8'hfc;
      17'd36826: data = 8'h01;
      17'd36827: data = 8'hfc;
      17'd36828: data = 8'hfc;
      17'd36829: data = 8'hfe;
      17'd36830: data = 8'hf9;
      17'd36831: data = 8'hfa;
      17'd36832: data = 8'h00;
      17'd36833: data = 8'hf9;
      17'd36834: data = 8'hf5;
      17'd36835: data = 8'hfa;
      17'd36836: data = 8'hfa;
      17'd36837: data = 8'hf9;
      17'd36838: data = 8'hfc;
      17'd36839: data = 8'hfd;
      17'd36840: data = 8'hfd;
      17'd36841: data = 8'h02;
      17'd36842: data = 8'h02;
      17'd36843: data = 8'h04;
      17'd36844: data = 8'h06;
      17'd36845: data = 8'h06;
      17'd36846: data = 8'h0c;
      17'd36847: data = 8'h06;
      17'd36848: data = 8'h02;
      17'd36849: data = 8'h05;
      17'd36850: data = 8'h06;
      17'd36851: data = 8'h04;
      17'd36852: data = 8'h01;
      17'd36853: data = 8'h01;
      17'd36854: data = 8'hfd;
      17'd36855: data = 8'hfd;
      17'd36856: data = 8'h02;
      17'd36857: data = 8'h01;
      17'd36858: data = 8'hfe;
      17'd36859: data = 8'hfd;
      17'd36860: data = 8'hfe;
      17'd36861: data = 8'h00;
      17'd36862: data = 8'hfe;
      17'd36863: data = 8'h00;
      17'd36864: data = 8'h00;
      17'd36865: data = 8'hfc;
      17'd36866: data = 8'hfd;
      17'd36867: data = 8'h01;
      17'd36868: data = 8'hfe;
      17'd36869: data = 8'hfc;
      17'd36870: data = 8'h00;
      17'd36871: data = 8'hfc;
      17'd36872: data = 8'hfc;
      17'd36873: data = 8'h00;
      17'd36874: data = 8'h00;
      17'd36875: data = 8'hfc;
      17'd36876: data = 8'hfc;
      17'd36877: data = 8'hfd;
      17'd36878: data = 8'hfd;
      17'd36879: data = 8'hfd;
      17'd36880: data = 8'hfc;
      17'd36881: data = 8'hf9;
      17'd36882: data = 8'hfc;
      17'd36883: data = 8'hf9;
      17'd36884: data = 8'hf4;
      17'd36885: data = 8'hf9;
      17'd36886: data = 8'hf6;
      17'd36887: data = 8'hfa;
      17'd36888: data = 8'hf9;
      17'd36889: data = 8'hf2;
      17'd36890: data = 8'hf4;
      17'd36891: data = 8'hf5;
      17'd36892: data = 8'hf4;
      17'd36893: data = 8'hf1;
      17'd36894: data = 8'hf1;
      17'd36895: data = 8'hf2;
      17'd36896: data = 8'hf5;
      17'd36897: data = 8'hf5;
      17'd36898: data = 8'hf4;
      17'd36899: data = 8'hfa;
      17'd36900: data = 8'h00;
      17'd36901: data = 8'hfc;
      17'd36902: data = 8'h00;
      17'd36903: data = 8'h0a;
      17'd36904: data = 8'h09;
      17'd36905: data = 8'h0a;
      17'd36906: data = 8'h0e;
      17'd36907: data = 8'h0d;
      17'd36908: data = 8'h11;
      17'd36909: data = 8'h1a;
      17'd36910: data = 8'h15;
      17'd36911: data = 8'h12;
      17'd36912: data = 8'h1a;
      17'd36913: data = 8'h16;
      17'd36914: data = 8'h16;
      17'd36915: data = 8'h16;
      17'd36916: data = 8'h13;
      17'd36917: data = 8'h19;
      17'd36918: data = 8'h15;
      17'd36919: data = 8'h13;
      17'd36920: data = 8'h13;
      17'd36921: data = 8'h0e;
      17'd36922: data = 8'h0e;
      17'd36923: data = 8'h12;
      17'd36924: data = 8'h0d;
      17'd36925: data = 8'h0c;
      17'd36926: data = 8'h0a;
      17'd36927: data = 8'h09;
      17'd36928: data = 8'h09;
      17'd36929: data = 8'h05;
      17'd36930: data = 8'h04;
      17'd36931: data = 8'h00;
      17'd36932: data = 8'hfe;
      17'd36933: data = 8'h01;
      17'd36934: data = 8'hf6;
      17'd36935: data = 8'hf9;
      17'd36936: data = 8'hfe;
      17'd36937: data = 8'hf4;
      17'd36938: data = 8'hfa;
      17'd36939: data = 8'hfc;
      17'd36940: data = 8'hf4;
      17'd36941: data = 8'hf6;
      17'd36942: data = 8'hf9;
      17'd36943: data = 8'hf2;
      17'd36944: data = 8'hf5;
      17'd36945: data = 8'hfc;
      17'd36946: data = 8'hf5;
      17'd36947: data = 8'hf2;
      17'd36948: data = 8'hf4;
      17'd36949: data = 8'hf2;
      17'd36950: data = 8'hf5;
      17'd36951: data = 8'hf4;
      17'd36952: data = 8'hef;
      17'd36953: data = 8'hf5;
      17'd36954: data = 8'hf5;
      17'd36955: data = 8'hf4;
      17'd36956: data = 8'hf9;
      17'd36957: data = 8'hf9;
      17'd36958: data = 8'hf6;
      17'd36959: data = 8'hf9;
      17'd36960: data = 8'hf6;
      17'd36961: data = 8'hf9;
      17'd36962: data = 8'hfa;
      17'd36963: data = 8'hf6;
      17'd36964: data = 8'hf6;
      17'd36965: data = 8'hfc;
      17'd36966: data = 8'hfc;
      17'd36967: data = 8'hf9;
      17'd36968: data = 8'hfc;
      17'd36969: data = 8'hfa;
      17'd36970: data = 8'hfa;
      17'd36971: data = 8'h00;
      17'd36972: data = 8'hfe;
      17'd36973: data = 8'hfc;
      17'd36974: data = 8'h01;
      17'd36975: data = 8'hfd;
      17'd36976: data = 8'hfc;
      17'd36977: data = 8'h04;
      17'd36978: data = 8'h01;
      17'd36979: data = 8'hfc;
      17'd36980: data = 8'hfd;
      17'd36981: data = 8'hfc;
      17'd36982: data = 8'hfd;
      17'd36983: data = 8'hfc;
      17'd36984: data = 8'hfc;
      17'd36985: data = 8'hf9;
      17'd36986: data = 8'hf5;
      17'd36987: data = 8'hf6;
      17'd36988: data = 8'hfa;
      17'd36989: data = 8'hfa;
      17'd36990: data = 8'hf2;
      17'd36991: data = 8'hf2;
      17'd36992: data = 8'hf1;
      17'd36993: data = 8'hf4;
      17'd36994: data = 8'hf9;
      17'd36995: data = 8'hf4;
      17'd36996: data = 8'hef;
      17'd36997: data = 8'hf2;
      17'd36998: data = 8'hf1;
      17'd36999: data = 8'hf6;
      17'd37000: data = 8'h05;
      17'd37001: data = 8'hfa;
      17'd37002: data = 8'hf1;
      17'd37003: data = 8'hfe;
      17'd37004: data = 8'hfe;
      17'd37005: data = 8'hf9;
      17'd37006: data = 8'h02;
      17'd37007: data = 8'h04;
      17'd37008: data = 8'hfc;
      17'd37009: data = 8'h04;
      17'd37010: data = 8'h00;
      17'd37011: data = 8'hfd;
      17'd37012: data = 8'h0c;
      17'd37013: data = 8'h0a;
      17'd37014: data = 8'h04;
      17'd37015: data = 8'h04;
      17'd37016: data = 8'h02;
      17'd37017: data = 8'h01;
      17'd37018: data = 8'h09;
      17'd37019: data = 8'h12;
      17'd37020: data = 8'h09;
      17'd37021: data = 8'hfc;
      17'd37022: data = 8'h05;
      17'd37023: data = 8'h09;
      17'd37024: data = 8'h04;
      17'd37025: data = 8'h06;
      17'd37026: data = 8'h00;
      17'd37027: data = 8'hfe;
      17'd37028: data = 8'h0a;
      17'd37029: data = 8'h0c;
      17'd37030: data = 8'h00;
      17'd37031: data = 8'hfa;
      17'd37032: data = 8'h02;
      17'd37033: data = 8'h02;
      17'd37034: data = 8'h01;
      17'd37035: data = 8'hf9;
      17'd37036: data = 8'hf4;
      17'd37037: data = 8'hf5;
      17'd37038: data = 8'hf4;
      17'd37039: data = 8'hf6;
      17'd37040: data = 8'hf6;
      17'd37041: data = 8'hed;
      17'd37042: data = 8'hef;
      17'd37043: data = 8'hfc;
      17'd37044: data = 8'hfe;
      17'd37045: data = 8'h00;
      17'd37046: data = 8'h02;
      17'd37047: data = 8'h09;
      17'd37048: data = 8'h0c;
      17'd37049: data = 8'h0d;
      17'd37050: data = 8'h11;
      17'd37051: data = 8'h0e;
      17'd37052: data = 8'h0e;
      17'd37053: data = 8'h0a;
      17'd37054: data = 8'h0a;
      17'd37055: data = 8'h0d;
      17'd37056: data = 8'h11;
      17'd37057: data = 8'h0e;
      17'd37058: data = 8'h0c;
      17'd37059: data = 8'h0a;
      17'd37060: data = 8'h09;
      17'd37061: data = 8'h0d;
      17'd37062: data = 8'h19;
      17'd37063: data = 8'h16;
      17'd37064: data = 8'h0e;
      17'd37065: data = 8'h15;
      17'd37066: data = 8'h13;
      17'd37067: data = 8'h13;
      17'd37068: data = 8'h13;
      17'd37069: data = 8'h09;
      17'd37070: data = 8'h05;
      17'd37071: data = 8'h02;
      17'd37072: data = 8'h05;
      17'd37073: data = 8'h05;
      17'd37074: data = 8'h00;
      17'd37075: data = 8'h02;
      17'd37076: data = 8'h00;
      17'd37077: data = 8'hfc;
      17'd37078: data = 8'hfc;
      17'd37079: data = 8'hfc;
      17'd37080: data = 8'hfd;
      17'd37081: data = 8'hfa;
      17'd37082: data = 8'hf4;
      17'd37083: data = 8'hf5;
      17'd37084: data = 8'hf4;
      17'd37085: data = 8'hf2;
      17'd37086: data = 8'hed;
      17'd37087: data = 8'he3;
      17'd37088: data = 8'he3;
      17'd37089: data = 8'he3;
      17'd37090: data = 8'he2;
      17'd37091: data = 8'he3;
      17'd37092: data = 8'hde;
      17'd37093: data = 8'hde;
      17'd37094: data = 8'he0;
      17'd37095: data = 8'he4;
      17'd37096: data = 8'he5;
      17'd37097: data = 8'he2;
      17'd37098: data = 8'hde;
      17'd37099: data = 8'he7;
      17'd37100: data = 8'hec;
      17'd37101: data = 8'hec;
      17'd37102: data = 8'hf1;
      17'd37103: data = 8'hf1;
      17'd37104: data = 8'hfa;
      17'd37105: data = 8'hfe;
      17'd37106: data = 8'hfe;
      17'd37107: data = 8'h02;
      17'd37108: data = 8'h09;
      17'd37109: data = 8'h13;
      17'd37110: data = 8'h19;
      17'd37111: data = 8'h1c;
      17'd37112: data = 8'h22;
      17'd37113: data = 8'h23;
      17'd37114: data = 8'h26;
      17'd37115: data = 8'h27;
      17'd37116: data = 8'h2b;
      17'd37117: data = 8'h2b;
      17'd37118: data = 8'h2c;
      17'd37119: data = 8'h2f;
      17'd37120: data = 8'h29;
      17'd37121: data = 8'h29;
      17'd37122: data = 8'h2f;
      17'd37123: data = 8'h29;
      17'd37124: data = 8'h22;
      17'd37125: data = 8'h23;
      17'd37126: data = 8'h1f;
      17'd37127: data = 8'h1a;
      17'd37128: data = 8'h1b;
      17'd37129: data = 8'h19;
      17'd37130: data = 8'h11;
      17'd37131: data = 8'h0d;
      17'd37132: data = 8'h0a;
      17'd37133: data = 8'h06;
      17'd37134: data = 8'h05;
      17'd37135: data = 8'hfd;
      17'd37136: data = 8'hf6;
      17'd37137: data = 8'hf6;
      17'd37138: data = 8'hf5;
      17'd37139: data = 8'hf2;
      17'd37140: data = 8'hf2;
      17'd37141: data = 8'hef;
      17'd37142: data = 8'he9;
      17'd37143: data = 8'heb;
      17'd37144: data = 8'he7;
      17'd37145: data = 8'he4;
      17'd37146: data = 8'he9;
      17'd37147: data = 8'he4;
      17'd37148: data = 8'he3;
      17'd37149: data = 8'he3;
      17'd37150: data = 8'he5;
      17'd37151: data = 8'he9;
      17'd37152: data = 8'he5;
      17'd37153: data = 8'he0;
      17'd37154: data = 8'he2;
      17'd37155: data = 8'he7;
      17'd37156: data = 8'hef;
      17'd37157: data = 8'hed;
      17'd37158: data = 8'hec;
      17'd37159: data = 8'hed;
      17'd37160: data = 8'hf1;
      17'd37161: data = 8'hf9;
      17'd37162: data = 8'hfd;
      17'd37163: data = 8'hfd;
      17'd37164: data = 8'hf9;
      17'd37165: data = 8'hf6;
      17'd37166: data = 8'h02;
      17'd37167: data = 8'h06;
      17'd37168: data = 8'h02;
      17'd37169: data = 8'h05;
      17'd37170: data = 8'h0c;
      17'd37171: data = 8'h06;
      17'd37172: data = 8'h0c;
      17'd37173: data = 8'h11;
      17'd37174: data = 8'h0d;
      17'd37175: data = 8'h0e;
      17'd37176: data = 8'h11;
      17'd37177: data = 8'h12;
      17'd37178: data = 8'h0c;
      17'd37179: data = 8'h06;
      17'd37180: data = 8'h0a;
      17'd37181: data = 8'h05;
      17'd37182: data = 8'h01;
      17'd37183: data = 8'hfe;
      17'd37184: data = 8'hfc;
      17'd37185: data = 8'hf9;
      17'd37186: data = 8'hf9;
      17'd37187: data = 8'hf9;
      17'd37188: data = 8'hf4;
      17'd37189: data = 8'hed;
      17'd37190: data = 8'hed;
      17'd37191: data = 8'hef;
      17'd37192: data = 8'he9;
      17'd37193: data = 8'he7;
      17'd37194: data = 8'he4;
      17'd37195: data = 8'he5;
      17'd37196: data = 8'he4;
      17'd37197: data = 8'hde;
      17'd37198: data = 8'he2;
      17'd37199: data = 8'hdc;
      17'd37200: data = 8'hdc;
      17'd37201: data = 8'he3;
      17'd37202: data = 8'he2;
      17'd37203: data = 8'he0;
      17'd37204: data = 8'hde;
      17'd37205: data = 8'he7;
      17'd37206: data = 8'heb;
      17'd37207: data = 8'heb;
      17'd37208: data = 8'hed;
      17'd37209: data = 8'hed;
      17'd37210: data = 8'hf1;
      17'd37211: data = 8'hf5;
      17'd37212: data = 8'hf6;
      17'd37213: data = 8'hfc;
      17'd37214: data = 8'hfe;
      17'd37215: data = 8'hfe;
      17'd37216: data = 8'hfe;
      17'd37217: data = 8'h04;
      17'd37218: data = 8'h04;
      17'd37219: data = 8'h04;
      17'd37220: data = 8'h0c;
      17'd37221: data = 8'h09;
      17'd37222: data = 8'h06;
      17'd37223: data = 8'h0a;
      17'd37224: data = 8'h06;
      17'd37225: data = 8'h06;
      17'd37226: data = 8'h09;
      17'd37227: data = 8'h06;
      17'd37228: data = 8'h06;
      17'd37229: data = 8'h0c;
      17'd37230: data = 8'h0a;
      17'd37231: data = 8'h09;
      17'd37232: data = 8'h0c;
      17'd37233: data = 8'h0d;
      17'd37234: data = 8'h0c;
      17'd37235: data = 8'h0d;
      17'd37236: data = 8'h0e;
      17'd37237: data = 8'h09;
      17'd37238: data = 8'h06;
      17'd37239: data = 8'h09;
      17'd37240: data = 8'h0d;
      17'd37241: data = 8'h04;
      17'd37242: data = 8'hfc;
      17'd37243: data = 8'h09;
      17'd37244: data = 8'h04;
      17'd37245: data = 8'h01;
      17'd37246: data = 8'h02;
      17'd37247: data = 8'hf9;
      17'd37248: data = 8'h01;
      17'd37249: data = 8'h02;
      17'd37250: data = 8'h01;
      17'd37251: data = 8'h02;
      17'd37252: data = 8'h00;
      17'd37253: data = 8'hfe;
      17'd37254: data = 8'h00;
      17'd37255: data = 8'hfe;
      17'd37256: data = 8'h06;
      17'd37257: data = 8'h04;
      17'd37258: data = 8'hfd;
      17'd37259: data = 8'h00;
      17'd37260: data = 8'h02;
      17'd37261: data = 8'h01;
      17'd37262: data = 8'h02;
      17'd37263: data = 8'h0e;
      17'd37264: data = 8'h06;
      17'd37265: data = 8'h01;
      17'd37266: data = 8'h06;
      17'd37267: data = 8'h01;
      17'd37268: data = 8'h01;
      17'd37269: data = 8'h0a;
      17'd37270: data = 8'h06;
      17'd37271: data = 8'h02;
      17'd37272: data = 8'h02;
      17'd37273: data = 8'h02;
      17'd37274: data = 8'h05;
      17'd37275: data = 8'h06;
      17'd37276: data = 8'h11;
      17'd37277: data = 8'h12;
      17'd37278: data = 8'h13;
      17'd37279: data = 8'h1b;
      17'd37280: data = 8'h19;
      17'd37281: data = 8'h1f;
      17'd37282: data = 8'h1f;
      17'd37283: data = 8'h1c;
      17'd37284: data = 8'h1e;
      17'd37285: data = 8'h1c;
      17'd37286: data = 8'h1c;
      17'd37287: data = 8'h19;
      17'd37288: data = 8'h19;
      17'd37289: data = 8'h1e;
      17'd37290: data = 8'h1e;
      17'd37291: data = 8'h1c;
      17'd37292: data = 8'h1a;
      17'd37293: data = 8'h16;
      17'd37294: data = 8'h1b;
      17'd37295: data = 8'h1b;
      17'd37296: data = 8'h1a;
      17'd37297: data = 8'h16;
      17'd37298: data = 8'h11;
      17'd37299: data = 8'h13;
      17'd37300: data = 8'h0d;
      17'd37301: data = 8'h0a;
      17'd37302: data = 8'h02;
      17'd37303: data = 8'hfa;
      17'd37304: data = 8'hfd;
      17'd37305: data = 8'hfc;
      17'd37306: data = 8'hf6;
      17'd37307: data = 8'hf4;
      17'd37308: data = 8'hed;
      17'd37309: data = 8'heb;
      17'd37310: data = 8'hed;
      17'd37311: data = 8'heb;
      17'd37312: data = 8'he4;
      17'd37313: data = 8'he3;
      17'd37314: data = 8'hde;
      17'd37315: data = 8'hdc;
      17'd37316: data = 8'hdc;
      17'd37317: data = 8'hda;
      17'd37318: data = 8'hd2;
      17'd37319: data = 8'hd8;
      17'd37320: data = 8'hd2;
      17'd37321: data = 8'hca;
      17'd37322: data = 8'hd2;
      17'd37323: data = 8'hd2;
      17'd37324: data = 8'hd8;
      17'd37325: data = 8'hdb;
      17'd37326: data = 8'hdb;
      17'd37327: data = 8'hde;
      17'd37328: data = 8'he5;
      17'd37329: data = 8'hed;
      17'd37330: data = 8'hed;
      17'd37331: data = 8'hf4;
      17'd37332: data = 8'hf6;
      17'd37333: data = 8'hf6;
      17'd37334: data = 8'h00;
      17'd37335: data = 8'h04;
      17'd37336: data = 8'h04;
      17'd37337: data = 8'h0a;
      17'd37338: data = 8'h0d;
      17'd37339: data = 8'h0e;
      17'd37340: data = 8'h19;
      17'd37341: data = 8'h1e;
      17'd37342: data = 8'h1f;
      17'd37343: data = 8'h27;
      17'd37344: data = 8'h2b;
      17'd37345: data = 8'h27;
      17'd37346: data = 8'h2f;
      17'd37347: data = 8'h34;
      17'd37348: data = 8'h31;
      17'd37349: data = 8'h2f;
      17'd37350: data = 8'h2f;
      17'd37351: data = 8'h2b;
      17'd37352: data = 8'h2c;
      17'd37353: data = 8'h2b;
      17'd37354: data = 8'h1f;
      17'd37355: data = 8'h22;
      17'd37356: data = 8'h23;
      17'd37357: data = 8'h1c;
      17'd37358: data = 8'h13;
      17'd37359: data = 8'h12;
      17'd37360: data = 8'h11;
      17'd37361: data = 8'h0a;
      17'd37362: data = 8'h05;
      17'd37363: data = 8'h04;
      17'd37364: data = 8'h00;
      17'd37365: data = 8'hfc;
      17'd37366: data = 8'hf6;
      17'd37367: data = 8'hf1;
      17'd37368: data = 8'hec;
      17'd37369: data = 8'hec;
      17'd37370: data = 8'heb;
      17'd37371: data = 8'he4;
      17'd37372: data = 8'he2;
      17'd37373: data = 8'he4;
      17'd37374: data = 8'hde;
      17'd37375: data = 8'hde;
      17'd37376: data = 8'he2;
      17'd37377: data = 8'hd8;
      17'd37378: data = 8'hda;
      17'd37379: data = 8'hde;
      17'd37380: data = 8'hdc;
      17'd37381: data = 8'hde;
      17'd37382: data = 8'he0;
      17'd37383: data = 8'hde;
      17'd37384: data = 8'he5;
      17'd37385: data = 8'hec;
      17'd37386: data = 8'he7;
      17'd37387: data = 8'hec;
      17'd37388: data = 8'hf1;
      17'd37389: data = 8'hf2;
      17'd37390: data = 8'hf9;
      17'd37391: data = 8'hfa;
      17'd37392: data = 8'hfa;
      17'd37393: data = 8'hfe;
      17'd37394: data = 8'h02;
      17'd37395: data = 8'h04;
      17'd37396: data = 8'h04;
      17'd37397: data = 8'h06;
      17'd37398: data = 8'h09;
      17'd37399: data = 8'h0c;
      17'd37400: data = 8'h0e;
      17'd37401: data = 8'h0a;
      17'd37402: data = 8'h0c;
      17'd37403: data = 8'h0e;
      17'd37404: data = 8'h0c;
      17'd37405: data = 8'h0c;
      17'd37406: data = 8'h0a;
      17'd37407: data = 8'h0a;
      17'd37408: data = 8'h0c;
      17'd37409: data = 8'h0c;
      17'd37410: data = 8'h05;
      17'd37411: data = 8'hfe;
      17'd37412: data = 8'hfe;
      17'd37413: data = 8'h00;
      17'd37414: data = 8'hfe;
      17'd37415: data = 8'hfc;
      17'd37416: data = 8'hfa;
      17'd37417: data = 8'hf4;
      17'd37418: data = 8'hef;
      17'd37419: data = 8'hf6;
      17'd37420: data = 8'hf4;
      17'd37421: data = 8'he5;
      17'd37422: data = 8'he2;
      17'd37423: data = 8'he5;
      17'd37424: data = 8'he3;
      17'd37425: data = 8'he7;
      17'd37426: data = 8'he4;
      17'd37427: data = 8'hdb;
      17'd37428: data = 8'he2;
      17'd37429: data = 8'he4;
      17'd37430: data = 8'hdc;
      17'd37431: data = 8'hde;
      17'd37432: data = 8'he7;
      17'd37433: data = 8'he3;
      17'd37434: data = 8'he4;
      17'd37435: data = 8'heb;
      17'd37436: data = 8'hed;
      17'd37437: data = 8'hef;
      17'd37438: data = 8'he9;
      17'd37439: data = 8'he9;
      17'd37440: data = 8'hf4;
      17'd37441: data = 8'hf5;
      17'd37442: data = 8'hf1;
      17'd37443: data = 8'hfa;
      17'd37444: data = 8'hfc;
      17'd37445: data = 8'hfc;
      17'd37446: data = 8'h06;
      17'd37447: data = 8'h06;
      17'd37448: data = 8'h02;
      17'd37449: data = 8'h06;
      17'd37450: data = 8'h0a;
      17'd37451: data = 8'h0e;
      17'd37452: data = 8'h13;
      17'd37453: data = 8'h0d;
      17'd37454: data = 8'h09;
      17'd37455: data = 8'h0e;
      17'd37456: data = 8'h11;
      17'd37457: data = 8'h0c;
      17'd37458: data = 8'h0a;
      17'd37459: data = 8'h05;
      17'd37460: data = 8'h05;
      17'd37461: data = 8'h09;
      17'd37462: data = 8'h09;
      17'd37463: data = 8'h05;
      17'd37464: data = 8'h05;
      17'd37465: data = 8'h05;
      17'd37466: data = 8'h02;
      17'd37467: data = 8'h01;
      17'd37468: data = 8'h00;
      17'd37469: data = 8'hfe;
      17'd37470: data = 8'hfe;
      17'd37471: data = 8'hfd;
      17'd37472: data = 8'h00;
      17'd37473: data = 8'h01;
      17'd37474: data = 8'hfd;
      17'd37475: data = 8'h00;
      17'd37476: data = 8'hfe;
      17'd37477: data = 8'hf9;
      17'd37478: data = 8'hfc;
      17'd37479: data = 8'hfd;
      17'd37480: data = 8'hfc;
      17'd37481: data = 8'h00;
      17'd37482: data = 8'h00;
      17'd37483: data = 8'hfe;
      17'd37484: data = 8'hfc;
      17'd37485: data = 8'hfd;
      17'd37486: data = 8'h00;
      17'd37487: data = 8'h02;
      17'd37488: data = 8'h06;
      17'd37489: data = 8'h01;
      17'd37490: data = 8'h05;
      17'd37491: data = 8'h13;
      17'd37492: data = 8'h0d;
      17'd37493: data = 8'h0e;
      17'd37494: data = 8'h0d;
      17'd37495: data = 8'h09;
      17'd37496: data = 8'h15;
      17'd37497: data = 8'h0e;
      17'd37498: data = 8'h0c;
      17'd37499: data = 8'h19;
      17'd37500: data = 8'h11;
      17'd37501: data = 8'h0c;
      17'd37502: data = 8'h1a;
      17'd37503: data = 8'h1b;
      17'd37504: data = 8'h0e;
      17'd37505: data = 8'h11;
      17'd37506: data = 8'h19;
      17'd37507: data = 8'h0d;
      17'd37508: data = 8'h12;
      17'd37509: data = 8'h1a;
      17'd37510: data = 8'h0c;
      17'd37511: data = 8'h11;
      17'd37512: data = 8'h15;
      17'd37513: data = 8'h0e;
      17'd37514: data = 8'h06;
      17'd37515: data = 8'h01;
      17'd37516: data = 8'h06;
      17'd37517: data = 8'h01;
      17'd37518: data = 8'hfa;
      17'd37519: data = 8'h01;
      17'd37520: data = 8'h04;
      17'd37521: data = 8'h00;
      17'd37522: data = 8'h04;
      17'd37523: data = 8'h06;
      17'd37524: data = 8'h05;
      17'd37525: data = 8'h04;
      17'd37526: data = 8'h06;
      17'd37527: data = 8'h0a;
      17'd37528: data = 8'h09;
      17'd37529: data = 8'h0c;
      17'd37530: data = 8'h09;
      17'd37531: data = 8'h09;
      17'd37532: data = 8'h0c;
      17'd37533: data = 8'h09;
      17'd37534: data = 8'h0a;
      17'd37535: data = 8'h04;
      17'd37536: data = 8'h02;
      17'd37537: data = 8'h0c;
      17'd37538: data = 8'h0d;
      17'd37539: data = 8'h0d;
      17'd37540: data = 8'h0e;
      17'd37541: data = 8'h0d;
      17'd37542: data = 8'h0a;
      17'd37543: data = 8'h0a;
      17'd37544: data = 8'h06;
      17'd37545: data = 8'h05;
      17'd37546: data = 8'h01;
      17'd37547: data = 8'h02;
      17'd37548: data = 8'h01;
      17'd37549: data = 8'h00;
      17'd37550: data = 8'h01;
      17'd37551: data = 8'hfc;
      17'd37552: data = 8'hfa;
      17'd37553: data = 8'hf9;
      17'd37554: data = 8'hf5;
      17'd37555: data = 8'hf4;
      17'd37556: data = 8'hef;
      17'd37557: data = 8'hed;
      17'd37558: data = 8'hed;
      17'd37559: data = 8'hec;
      17'd37560: data = 8'heb;
      17'd37561: data = 8'he5;
      17'd37562: data = 8'he2;
      17'd37563: data = 8'he2;
      17'd37564: data = 8'he0;
      17'd37565: data = 8'hdc;
      17'd37566: data = 8'he0;
      17'd37567: data = 8'he0;
      17'd37568: data = 8'he0;
      17'd37569: data = 8'he2;
      17'd37570: data = 8'he4;
      17'd37571: data = 8'he5;
      17'd37572: data = 8'he5;
      17'd37573: data = 8'he7;
      17'd37574: data = 8'hec;
      17'd37575: data = 8'hed;
      17'd37576: data = 8'hf2;
      17'd37577: data = 8'hfa;
      17'd37578: data = 8'hfa;
      17'd37579: data = 8'hfc;
      17'd37580: data = 8'hfd;
      17'd37581: data = 8'hfe;
      17'd37582: data = 8'h04;
      17'd37583: data = 8'h05;
      17'd37584: data = 8'h09;
      17'd37585: data = 8'h0d;
      17'd37586: data = 8'h12;
      17'd37587: data = 8'h1a;
      17'd37588: data = 8'h1c;
      17'd37589: data = 8'h1b;
      17'd37590: data = 8'h22;
      17'd37591: data = 8'h23;
      17'd37592: data = 8'h23;
      17'd37593: data = 8'h24;
      17'd37594: data = 8'h23;
      17'd37595: data = 8'h23;
      17'd37596: data = 8'h24;
      17'd37597: data = 8'h22;
      17'd37598: data = 8'h1c;
      17'd37599: data = 8'h1c;
      17'd37600: data = 8'h1a;
      17'd37601: data = 8'h13;
      17'd37602: data = 8'h12;
      17'd37603: data = 8'h11;
      17'd37604: data = 8'h0e;
      17'd37605: data = 8'h0d;
      17'd37606: data = 8'h0a;
      17'd37607: data = 8'h09;
      17'd37608: data = 8'h05;
      17'd37609: data = 8'h02;
      17'd37610: data = 8'hfe;
      17'd37611: data = 8'hfc;
      17'd37612: data = 8'hfc;
      17'd37613: data = 8'hf6;
      17'd37614: data = 8'hed;
      17'd37615: data = 8'hed;
      17'd37616: data = 8'hec;
      17'd37617: data = 8'he9;
      17'd37618: data = 8'he5;
      17'd37619: data = 8'he0;
      17'd37620: data = 8'he0;
      17'd37621: data = 8'hde;
      17'd37622: data = 8'he3;
      17'd37623: data = 8'he3;
      17'd37624: data = 8'he3;
      17'd37625: data = 8'he5;
      17'd37626: data = 8'he5;
      17'd37627: data = 8'he5;
      17'd37628: data = 8'he7;
      17'd37629: data = 8'he9;
      17'd37630: data = 8'he7;
      17'd37631: data = 8'hec;
      17'd37632: data = 8'hed;
      17'd37633: data = 8'hf1;
      17'd37634: data = 8'hf1;
      17'd37635: data = 8'hf1;
      17'd37636: data = 8'hf9;
      17'd37637: data = 8'hfe;
      17'd37638: data = 8'hfd;
      17'd37639: data = 8'hfc;
      17'd37640: data = 8'h00;
      17'd37641: data = 8'h06;
      17'd37642: data = 8'h09;
      17'd37643: data = 8'h0d;
      17'd37644: data = 8'h11;
      17'd37645: data = 8'h0c;
      17'd37646: data = 8'h11;
      17'd37647: data = 8'h15;
      17'd37648: data = 8'h11;
      17'd37649: data = 8'h12;
      17'd37650: data = 8'h12;
      17'd37651: data = 8'h0c;
      17'd37652: data = 8'h0c;
      17'd37653: data = 8'h0d;
      17'd37654: data = 8'h0c;
      17'd37655: data = 8'h09;
      17'd37656: data = 8'h09;
      17'd37657: data = 8'hfc;
      17'd37658: data = 8'hf5;
      17'd37659: data = 8'hfe;
      17'd37660: data = 8'hfc;
      17'd37661: data = 8'hfa;
      17'd37662: data = 8'hfe;
      17'd37663: data = 8'hfc;
      17'd37664: data = 8'hed;
      17'd37665: data = 8'hf1;
      17'd37666: data = 8'hfa;
      17'd37667: data = 8'hf4;
      17'd37668: data = 8'he7;
      17'd37669: data = 8'he7;
      17'd37670: data = 8'he5;
      17'd37671: data = 8'he7;
      17'd37672: data = 8'heb;
      17'd37673: data = 8'he7;
      17'd37674: data = 8'hde;
      17'd37675: data = 8'hde;
      17'd37676: data = 8'he9;
      17'd37677: data = 8'he4;
      17'd37678: data = 8'he3;
      17'd37679: data = 8'hec;
      17'd37680: data = 8'hed;
      17'd37681: data = 8'heb;
      17'd37682: data = 8'hf5;
      17'd37683: data = 8'hfe;
      17'd37684: data = 8'hf4;
      17'd37685: data = 8'hef;
      17'd37686: data = 8'hf9;
      17'd37687: data = 8'hfd;
      17'd37688: data = 8'hfc;
      17'd37689: data = 8'h00;
      17'd37690: data = 8'h00;
      17'd37691: data = 8'h04;
      17'd37692: data = 8'h09;
      17'd37693: data = 8'h09;
      17'd37694: data = 8'h06;
      17'd37695: data = 8'h05;
      17'd37696: data = 8'h09;
      17'd37697: data = 8'h09;
      17'd37698: data = 8'h09;
      17'd37699: data = 8'h0c;
      17'd37700: data = 8'h0a;
      17'd37701: data = 8'h05;
      17'd37702: data = 8'h06;
      17'd37703: data = 8'h05;
      17'd37704: data = 8'h05;
      17'd37705: data = 8'h04;
      17'd37706: data = 8'h02;
      17'd37707: data = 8'h00;
      17'd37708: data = 8'h02;
      17'd37709: data = 8'h0a;
      17'd37710: data = 8'h05;
      17'd37711: data = 8'h02;
      17'd37712: data = 8'h01;
      17'd37713: data = 8'hfc;
      17'd37714: data = 8'hfc;
      17'd37715: data = 8'h00;
      17'd37716: data = 8'hfe;
      17'd37717: data = 8'hfc;
      17'd37718: data = 8'hf6;
      17'd37719: data = 8'hf4;
      17'd37720: data = 8'hfc;
      17'd37721: data = 8'hfd;
      17'd37722: data = 8'hf6;
      17'd37723: data = 8'hf6;
      17'd37724: data = 8'hf2;
      17'd37725: data = 8'hf6;
      17'd37726: data = 8'h01;
      17'd37727: data = 8'hfc;
      17'd37728: data = 8'hf9;
      17'd37729: data = 8'hfd;
      17'd37730: data = 8'hfd;
      17'd37731: data = 8'hfc;
      17'd37732: data = 8'h01;
      17'd37733: data = 8'h00;
      17'd37734: data = 8'hfd;
      17'd37735: data = 8'h00;
      17'd37736: data = 8'h02;
      17'd37737: data = 8'h0a;
      17'd37738: data = 8'h05;
      17'd37739: data = 8'h02;
      17'd37740: data = 8'h06;
      17'd37741: data = 8'h06;
      17'd37742: data = 8'h0e;
      17'd37743: data = 8'h0c;
      17'd37744: data = 8'h0c;
      17'd37745: data = 8'h15;
      17'd37746: data = 8'h0c;
      17'd37747: data = 8'h11;
      17'd37748: data = 8'h15;
      17'd37749: data = 8'h0e;
      17'd37750: data = 8'h0e;
      17'd37751: data = 8'h06;
      17'd37752: data = 8'h0d;
      17'd37753: data = 8'h12;
      17'd37754: data = 8'h0c;
      17'd37755: data = 8'h19;
      17'd37756: data = 8'h11;
      17'd37757: data = 8'h05;
      17'd37758: data = 8'h0d;
      17'd37759: data = 8'h0e;
      17'd37760: data = 8'h0a;
      17'd37761: data = 8'h05;
      17'd37762: data = 8'h0c;
      17'd37763: data = 8'h0c;
      17'd37764: data = 8'h00;
      17'd37765: data = 8'h09;
      17'd37766: data = 8'h06;
      17'd37767: data = 8'hfc;
      17'd37768: data = 8'h02;
      17'd37769: data = 8'h00;
      17'd37770: data = 8'hfd;
      17'd37771: data = 8'hf1;
      17'd37772: data = 8'hf9;
      17'd37773: data = 8'h06;
      17'd37774: data = 8'hf1;
      17'd37775: data = 8'hfd;
      17'd37776: data = 8'h05;
      17'd37777: data = 8'hf5;
      17'd37778: data = 8'hfe;
      17'd37779: data = 8'h05;
      17'd37780: data = 8'h06;
      17'd37781: data = 8'h00;
      17'd37782: data = 8'h05;
      17'd37783: data = 8'h13;
      17'd37784: data = 8'h00;
      17'd37785: data = 8'h02;
      17'd37786: data = 8'h0c;
      17'd37787: data = 8'hfd;
      17'd37788: data = 8'h04;
      17'd37789: data = 8'h06;
      17'd37790: data = 8'h0a;
      17'd37791: data = 8'h05;
      17'd37792: data = 8'h02;
      17'd37793: data = 8'h11;
      17'd37794: data = 8'h0d;
      17'd37795: data = 8'h0a;
      17'd37796: data = 8'h11;
      17'd37797: data = 8'h0a;
      17'd37798: data = 8'h11;
      17'd37799: data = 8'h0c;
      17'd37800: data = 8'h09;
      17'd37801: data = 8'h0c;
      17'd37802: data = 8'h05;
      17'd37803: data = 8'h09;
      17'd37804: data = 8'h00;
      17'd37805: data = 8'hfc;
      17'd37806: data = 8'h00;
      17'd37807: data = 8'hf5;
      17'd37808: data = 8'hf9;
      17'd37809: data = 8'hfc;
      17'd37810: data = 8'hf6;
      17'd37811: data = 8'hfa;
      17'd37812: data = 8'hf2;
      17'd37813: data = 8'hf1;
      17'd37814: data = 8'hf2;
      17'd37815: data = 8'heb;
      17'd37816: data = 8'hed;
      17'd37817: data = 8'he9;
      17'd37818: data = 8'he9;
      17'd37819: data = 8'he9;
      17'd37820: data = 8'he0;
      17'd37821: data = 8'he5;
      17'd37822: data = 8'he2;
      17'd37823: data = 8'he4;
      17'd37824: data = 8'he5;
      17'd37825: data = 8'hde;
      17'd37826: data = 8'he5;
      17'd37827: data = 8'he4;
      17'd37828: data = 8'he9;
      17'd37829: data = 8'hf5;
      17'd37830: data = 8'heb;
      17'd37831: data = 8'he9;
      17'd37832: data = 8'hf4;
      17'd37833: data = 8'hf9;
      17'd37834: data = 8'hf5;
      17'd37835: data = 8'hf5;
      17'd37836: data = 8'hfd;
      17'd37837: data = 8'hfa;
      17'd37838: data = 8'h00;
      17'd37839: data = 8'h0c;
      17'd37840: data = 8'h04;
      17'd37841: data = 8'h04;
      17'd37842: data = 8'h0d;
      17'd37843: data = 8'h12;
      17'd37844: data = 8'h1b;
      17'd37845: data = 8'h16;
      17'd37846: data = 8'h19;
      17'd37847: data = 8'h1b;
      17'd37848: data = 8'h1a;
      17'd37849: data = 8'h24;
      17'd37850: data = 8'h22;
      17'd37851: data = 8'h1b;
      17'd37852: data = 8'h1b;
      17'd37853: data = 8'h19;
      17'd37854: data = 8'h1c;
      17'd37855: data = 8'h16;
      17'd37856: data = 8'h16;
      17'd37857: data = 8'h15;
      17'd37858: data = 8'h0e;
      17'd37859: data = 8'h13;
      17'd37860: data = 8'h0d;
      17'd37861: data = 8'h09;
      17'd37862: data = 8'h09;
      17'd37863: data = 8'h02;
      17'd37864: data = 8'h01;
      17'd37865: data = 8'hfe;
      17'd37866: data = 8'hfd;
      17'd37867: data = 8'hfc;
      17'd37868: data = 8'hf5;
      17'd37869: data = 8'hf2;
      17'd37870: data = 8'hf1;
      17'd37871: data = 8'hf2;
      17'd37872: data = 8'hed;
      17'd37873: data = 8'he9;
      17'd37874: data = 8'he9;
      17'd37875: data = 8'he9;
      17'd37876: data = 8'he9;
      17'd37877: data = 8'heb;
      17'd37878: data = 8'he7;
      17'd37879: data = 8'he9;
      17'd37880: data = 8'he7;
      17'd37881: data = 8'he7;
      17'd37882: data = 8'hec;
      17'd37883: data = 8'hed;
      17'd37884: data = 8'hef;
      17'd37885: data = 8'hed;
      17'd37886: data = 8'hed;
      17'd37887: data = 8'hf2;
      17'd37888: data = 8'hf4;
      17'd37889: data = 8'hfa;
      17'd37890: data = 8'hfa;
      17'd37891: data = 8'hf4;
      17'd37892: data = 8'hfd;
      17'd37893: data = 8'h00;
      17'd37894: data = 8'h01;
      17'd37895: data = 8'h01;
      17'd37896: data = 8'hfe;
      17'd37897: data = 8'h04;
      17'd37898: data = 8'h06;
      17'd37899: data = 8'h09;
      17'd37900: data = 8'h06;
      17'd37901: data = 8'h06;
      17'd37902: data = 8'h0a;
      17'd37903: data = 8'h09;
      17'd37904: data = 8'h0a;
      17'd37905: data = 8'h09;
      17'd37906: data = 8'h09;
      17'd37907: data = 8'h06;
      17'd37908: data = 8'h06;
      17'd37909: data = 8'h0c;
      17'd37910: data = 8'h04;
      17'd37911: data = 8'hfa;
      17'd37912: data = 8'hfe;
      17'd37913: data = 8'h02;
      17'd37914: data = 8'h02;
      17'd37915: data = 8'h01;
      17'd37916: data = 8'hfc;
      17'd37917: data = 8'hfd;
      17'd37918: data = 8'hfd;
      17'd37919: data = 8'hfd;
      17'd37920: data = 8'hfc;
      17'd37921: data = 8'hf9;
      17'd37922: data = 8'hf2;
      17'd37923: data = 8'hf2;
      17'd37924: data = 8'hf4;
      17'd37925: data = 8'hf1;
      17'd37926: data = 8'hed;
      17'd37927: data = 8'he9;
      17'd37928: data = 8'he4;
      17'd37929: data = 8'he9;
      17'd37930: data = 8'heb;
      17'd37931: data = 8'he4;
      17'd37932: data = 8'he4;
      17'd37933: data = 8'heb;
      17'd37934: data = 8'heb;
      17'd37935: data = 8'heb;
      17'd37936: data = 8'he9;
      17'd37937: data = 8'heb;
      17'd37938: data = 8'he7;
      17'd37939: data = 8'he7;
      17'd37940: data = 8'hed;
      17'd37941: data = 8'hf1;
      17'd37942: data = 8'hf1;
      17'd37943: data = 8'hf2;
      17'd37944: data = 8'hf4;
      17'd37945: data = 8'hfa;
      17'd37946: data = 8'hfe;
      17'd37947: data = 8'hfe;
      17'd37948: data = 8'hfe;
      17'd37949: data = 8'h00;
      17'd37950: data = 8'h02;
      17'd37951: data = 8'h04;
      17'd37952: data = 8'h06;
      17'd37953: data = 8'h05;
      17'd37954: data = 8'h02;
      17'd37955: data = 8'h02;
      17'd37956: data = 8'h01;
      17'd37957: data = 8'h00;
      17'd37958: data = 8'h00;
      17'd37959: data = 8'h00;
      17'd37960: data = 8'h02;
      17'd37961: data = 8'h04;
      17'd37962: data = 8'h02;
      17'd37963: data = 8'h04;
      17'd37964: data = 8'h01;
      17'd37965: data = 8'h04;
      17'd37966: data = 8'h04;
      17'd37967: data = 8'hfd;
      17'd37968: data = 8'hfe;
      17'd37969: data = 8'hfe;
      17'd37970: data = 8'h00;
      17'd37971: data = 8'hfd;
      17'd37972: data = 8'hfc;
      17'd37973: data = 8'hfa;
      17'd37974: data = 8'hfa;
      17'd37975: data = 8'hfa;
      17'd37976: data = 8'hf6;
      17'd37977: data = 8'hf6;
      17'd37978: data = 8'hfd;
      17'd37979: data = 8'h09;
      17'd37980: data = 8'h09;
      17'd37981: data = 8'hfe;
      17'd37982: data = 8'hfa;
      17'd37983: data = 8'hfd;
      17'd37984: data = 8'h06;
      17'd37985: data = 8'h19;
      17'd37986: data = 8'h04;
      17'd37987: data = 8'hf1;
      17'd37988: data = 8'h01;
      17'd37989: data = 8'h0d;
      17'd37990: data = 8'h0c;
      17'd37991: data = 8'h0c;
      17'd37992: data = 8'h09;
      17'd37993: data = 8'hf9;
      17'd37994: data = 8'hfa;
      17'd37995: data = 8'h15;
      17'd37996: data = 8'h19;
      17'd37997: data = 8'h05;
      17'd37998: data = 8'hf1;
      17'd37999: data = 8'hfd;
      17'd38000: data = 8'h23;
      17'd38001: data = 8'h31;
      17'd38002: data = 8'h01;
      17'd38003: data = 8'hdb;
      17'd38004: data = 8'h0d;
      17'd38005: data = 8'h33;
      17'd38006: data = 8'h23;
      17'd38007: data = 8'h1e;
      17'd38008: data = 8'hfd;
      17'd38009: data = 8'hf2;
      17'd38010: data = 8'h2b;
      17'd38011: data = 8'h1e;
      17'd38012: data = 8'h0c;
      17'd38013: data = 8'h0d;
      17'd38014: data = 8'h09;
      17'd38015: data = 8'h1e;
      17'd38016: data = 8'h15;
      17'd38017: data = 8'h05;
      17'd38018: data = 8'h06;
      17'd38019: data = 8'h1b;
      17'd38020: data = 8'h1f;
      17'd38021: data = 8'h0c;
      17'd38022: data = 8'h00;
      17'd38023: data = 8'hfc;
      17'd38024: data = 8'h0d;
      17'd38025: data = 8'h1f;
      17'd38026: data = 8'h12;
      17'd38027: data = 8'hfe;
      17'd38028: data = 8'hfd;
      17'd38029: data = 8'h01;
      17'd38030: data = 8'h09;
      17'd38031: data = 8'h04;
      17'd38032: data = 8'hfe;
      17'd38033: data = 8'hfd;
      17'd38034: data = 8'h00;
      17'd38035: data = 8'h0a;
      17'd38036: data = 8'h05;
      17'd38037: data = 8'hf9;
      17'd38038: data = 8'hf1;
      17'd38039: data = 8'h01;
      17'd38040: data = 8'h06;
      17'd38041: data = 8'hf5;
      17'd38042: data = 8'hec;
      17'd38043: data = 8'hf9;
      17'd38044: data = 8'h04;
      17'd38045: data = 8'h04;
      17'd38046: data = 8'hfa;
      17'd38047: data = 8'hf9;
      17'd38048: data = 8'h05;
      17'd38049: data = 8'h04;
      17'd38050: data = 8'h04;
      17'd38051: data = 8'h06;
      17'd38052: data = 8'h01;
      17'd38053: data = 8'h06;
      17'd38054: data = 8'h0e;
      17'd38055: data = 8'h0c;
      17'd38056: data = 8'h02;
      17'd38057: data = 8'h06;
      17'd38058: data = 8'h0d;
      17'd38059: data = 8'h02;
      17'd38060: data = 8'h00;
      17'd38061: data = 8'h0a;
      17'd38062: data = 8'h0c;
      17'd38063: data = 8'h06;
      17'd38064: data = 8'h09;
      17'd38065: data = 8'h0a;
      17'd38066: data = 8'h04;
      17'd38067: data = 8'h04;
      17'd38068: data = 8'h0e;
      17'd38069: data = 8'h09;
      17'd38070: data = 8'hfd;
      17'd38071: data = 8'hfe;
      17'd38072: data = 8'h00;
      17'd38073: data = 8'hfe;
      17'd38074: data = 8'hfd;
      17'd38075: data = 8'h00;
      17'd38076: data = 8'hfc;
      17'd38077: data = 8'hf1;
      17'd38078: data = 8'hf2;
      17'd38079: data = 8'hfa;
      17'd38080: data = 8'hfc;
      17'd38081: data = 8'hf5;
      17'd38082: data = 8'hf2;
      17'd38083: data = 8'hf1;
      17'd38084: data = 8'hef;
      17'd38085: data = 8'hf1;
      17'd38086: data = 8'hf4;
      17'd38087: data = 8'he9;
      17'd38088: data = 8'hde;
      17'd38089: data = 8'he0;
      17'd38090: data = 8'he4;
      17'd38091: data = 8'he7;
      17'd38092: data = 8'he3;
      17'd38093: data = 8'hde;
      17'd38094: data = 8'hda;
      17'd38095: data = 8'hde;
      17'd38096: data = 8'he4;
      17'd38097: data = 8'he5;
      17'd38098: data = 8'he4;
      17'd38099: data = 8'he2;
      17'd38100: data = 8'he5;
      17'd38101: data = 8'hed;
      17'd38102: data = 8'hf2;
      17'd38103: data = 8'hf1;
      17'd38104: data = 8'hf1;
      17'd38105: data = 8'hf5;
      17'd38106: data = 8'hf9;
      17'd38107: data = 8'hfd;
      17'd38108: data = 8'h01;
      17'd38109: data = 8'h00;
      17'd38110: data = 8'h01;
      17'd38111: data = 8'h09;
      17'd38112: data = 8'h0c;
      17'd38113: data = 8'h09;
      17'd38114: data = 8'h0d;
      17'd38115: data = 8'h0d;
      17'd38116: data = 8'h0c;
      17'd38117: data = 8'h11;
      17'd38118: data = 8'h13;
      17'd38119: data = 8'h11;
      17'd38120: data = 8'h0e;
      17'd38121: data = 8'h12;
      17'd38122: data = 8'h15;
      17'd38123: data = 8'h13;
      17'd38124: data = 8'h15;
      17'd38125: data = 8'h11;
      17'd38126: data = 8'h0e;
      17'd38127: data = 8'h11;
      17'd38128: data = 8'h0e;
      17'd38129: data = 8'h0e;
      17'd38130: data = 8'h0c;
      17'd38131: data = 8'h09;
      17'd38132: data = 8'h04;
      17'd38133: data = 8'h02;
      17'd38134: data = 8'h01;
      17'd38135: data = 8'h01;
      17'd38136: data = 8'h00;
      17'd38137: data = 8'hfc;
      17'd38138: data = 8'hfa;
      17'd38139: data = 8'hf6;
      17'd38140: data = 8'hf6;
      17'd38141: data = 8'hfd;
      17'd38142: data = 8'hfa;
      17'd38143: data = 8'hf1;
      17'd38144: data = 8'hf1;
      17'd38145: data = 8'hf6;
      17'd38146: data = 8'hf6;
      17'd38147: data = 8'hf5;
      17'd38148: data = 8'hf2;
      17'd38149: data = 8'he9;
      17'd38150: data = 8'he9;
      17'd38151: data = 8'hf2;
      17'd38152: data = 8'hf4;
      17'd38153: data = 8'hf1;
      17'd38154: data = 8'hed;
      17'd38155: data = 8'hf1;
      17'd38156: data = 8'hf2;
      17'd38157: data = 8'hf5;
      17'd38158: data = 8'hfa;
      17'd38159: data = 8'hf9;
      17'd38160: data = 8'hf5;
      17'd38161: data = 8'hf6;
      17'd38162: data = 8'hfc;
      17'd38163: data = 8'hfd;
      17'd38164: data = 8'hfd;
      17'd38165: data = 8'hfc;
      17'd38166: data = 8'hfa;
      17'd38167: data = 8'hfe;
      17'd38168: data = 8'h04;
      17'd38169: data = 8'h01;
      17'd38170: data = 8'hfd;
      17'd38171: data = 8'hfe;
      17'd38172: data = 8'hfd;
      17'd38173: data = 8'hfe;
      17'd38174: data = 8'h01;
      17'd38175: data = 8'h00;
      17'd38176: data = 8'hfe;
      17'd38177: data = 8'h01;
      17'd38178: data = 8'h02;
      17'd38179: data = 8'hfc;
      17'd38180: data = 8'h00;
      17'd38181: data = 8'h06;
      17'd38182: data = 8'h04;
      17'd38183: data = 8'hfc;
      17'd38184: data = 8'hfa;
      17'd38185: data = 8'hfd;
      17'd38186: data = 8'hfd;
      17'd38187: data = 8'h00;
      17'd38188: data = 8'hfc;
      17'd38189: data = 8'hf5;
      17'd38190: data = 8'hf9;
      17'd38191: data = 8'hfc;
      17'd38192: data = 8'hf9;
      17'd38193: data = 8'hf5;
      17'd38194: data = 8'hf5;
      17'd38195: data = 8'hf4;
      17'd38196: data = 8'hf6;
      17'd38197: data = 8'hf6;
      17'd38198: data = 8'hf4;
      17'd38199: data = 8'hef;
      17'd38200: data = 8'hf1;
      17'd38201: data = 8'hf6;
      17'd38202: data = 8'hf4;
      17'd38203: data = 8'hf1;
      17'd38204: data = 8'hf5;
      17'd38205: data = 8'hef;
      17'd38206: data = 8'hf5;
      17'd38207: data = 8'h00;
      17'd38208: data = 8'hf6;
      17'd38209: data = 8'hf6;
      17'd38210: data = 8'hf9;
      17'd38211: data = 8'hf4;
      17'd38212: data = 8'hfc;
      17'd38213: data = 8'h05;
      17'd38214: data = 8'hfe;
      17'd38215: data = 8'hf5;
      17'd38216: data = 8'hfa;
      17'd38217: data = 8'hfe;
      17'd38218: data = 8'hfa;
      17'd38219: data = 8'hf4;
      17'd38220: data = 8'hf9;
      17'd38221: data = 8'h1a;
      17'd38222: data = 8'h1f;
      17'd38223: data = 8'he3;
      17'd38224: data = 8'he3;
      17'd38225: data = 8'h19;
      17'd38226: data = 8'h15;
      17'd38227: data = 8'h05;
      17'd38228: data = 8'h00;
      17'd38229: data = 8'hfe;
      17'd38230: data = 8'h09;
      17'd38231: data = 8'hfd;
      17'd38232: data = 8'h16;
      17'd38233: data = 8'h26;
      17'd38234: data = 8'he7;
      17'd38235: data = 8'h09;
      17'd38236: data = 8'h0e;
      17'd38237: data = 8'hf4;
      17'd38238: data = 8'h24;
      17'd38239: data = 8'h29;
      17'd38240: data = 8'h05;
      17'd38241: data = 8'heb;
      17'd38242: data = 8'h00;
      17'd38243: data = 8'h13;
      17'd38244: data = 8'h19;
      17'd38245: data = 8'h2d;
      17'd38246: data = 8'hfe;
      17'd38247: data = 8'hdb;
      17'd38248: data = 8'h19;
      17'd38249: data = 8'h13;
      17'd38250: data = 8'h0c;
      17'd38251: data = 8'h2c;
      17'd38252: data = 8'h01;
      17'd38253: data = 8'hfd;
      17'd38254: data = 8'hfe;
      17'd38255: data = 8'hf1;
      17'd38256: data = 8'h1b;
      17'd38257: data = 8'h26;
      17'd38258: data = 8'hf4;
      17'd38259: data = 8'h0c;
      17'd38260: data = 8'h1f;
      17'd38261: data = 8'he4;
      17'd38262: data = 8'heb;
      17'd38263: data = 8'h1a;
      17'd38264: data = 8'h24;
      17'd38265: data = 8'h0e;
      17'd38266: data = 8'hfa;
      17'd38267: data = 8'hf4;
      17'd38268: data = 8'h12;
      17'd38269: data = 8'h1f;
      17'd38270: data = 8'h16;
      17'd38271: data = 8'h06;
      17'd38272: data = 8'hfd;
      17'd38273: data = 8'h11;
      17'd38274: data = 8'h01;
      17'd38275: data = 8'h01;
      17'd38276: data = 8'h24;
      17'd38277: data = 8'h24;
      17'd38278: data = 8'h01;
      17'd38279: data = 8'hef;
      17'd38280: data = 8'h11;
      17'd38281: data = 8'h12;
      17'd38282: data = 8'h13;
      17'd38283: data = 8'h15;
      17'd38284: data = 8'h0c;
      17'd38285: data = 8'he5;
      17'd38286: data = 8'h00;
      17'd38287: data = 8'h42;
      17'd38288: data = 8'h13;
      17'd38289: data = 8'hf6;
      17'd38290: data = 8'hfd;
      17'd38291: data = 8'hf4;
      17'd38292: data = 8'h00;
      17'd38293: data = 8'h1c;
      17'd38294: data = 8'h0d;
      17'd38295: data = 8'h04;
      17'd38296: data = 8'hf2;
      17'd38297: data = 8'hf6;
      17'd38298: data = 8'h19;
      17'd38299: data = 8'h12;
      17'd38300: data = 8'hfc;
      17'd38301: data = 8'hf6;
      17'd38302: data = 8'h11;
      17'd38303: data = 8'hfa;
      17'd38304: data = 8'he5;
      17'd38305: data = 8'h0c;
      17'd38306: data = 8'h1a;
      17'd38307: data = 8'h05;
      17'd38308: data = 8'hf5;
      17'd38309: data = 8'hf2;
      17'd38310: data = 8'hed;
      17'd38311: data = 8'h0c;
      17'd38312: data = 8'h12;
      17'd38313: data = 8'hf4;
      17'd38314: data = 8'hfe;
      17'd38315: data = 8'hfa;
      17'd38316: data = 8'hf4;
      17'd38317: data = 8'h23;
      17'd38318: data = 8'h06;
      17'd38319: data = 8'hd8;
      17'd38320: data = 8'h05;
      17'd38321: data = 8'hfe;
      17'd38322: data = 8'hf5;
      17'd38323: data = 8'h05;
      17'd38324: data = 8'hf9;
      17'd38325: data = 8'hfe;
      17'd38326: data = 8'h04;
      17'd38327: data = 8'h00;
      17'd38328: data = 8'hf4;
      17'd38329: data = 8'hef;
      17'd38330: data = 8'hfd;
      17'd38331: data = 8'h04;
      17'd38332: data = 8'hf6;
      17'd38333: data = 8'hf2;
      17'd38334: data = 8'hfa;
      17'd38335: data = 8'hf9;
      17'd38336: data = 8'h01;
      17'd38337: data = 8'h02;
      17'd38338: data = 8'he7;
      17'd38339: data = 8'hde;
      17'd38340: data = 8'hfa;
      17'd38341: data = 8'h01;
      17'd38342: data = 8'hfd;
      17'd38343: data = 8'hf4;
      17'd38344: data = 8'hf2;
      17'd38345: data = 8'h06;
      17'd38346: data = 8'hfe;
      17'd38347: data = 8'heb;
      17'd38348: data = 8'hfc;
      17'd38349: data = 8'h01;
      17'd38350: data = 8'hf9;
      17'd38351: data = 8'hf6;
      17'd38352: data = 8'hf1;
      17'd38353: data = 8'hf6;
      17'd38354: data = 8'h04;
      17'd38355: data = 8'h09;
      17'd38356: data = 8'hfa;
      17'd38357: data = 8'he2;
      17'd38358: data = 8'he7;
      17'd38359: data = 8'h01;
      17'd38360: data = 8'h0c;
      17'd38361: data = 8'hf9;
      17'd38362: data = 8'hef;
      17'd38363: data = 8'hf6;
      17'd38364: data = 8'hf9;
      17'd38365: data = 8'h01;
      17'd38366: data = 8'h04;
      17'd38367: data = 8'hf5;
      17'd38368: data = 8'he9;
      17'd38369: data = 8'hef;
      17'd38370: data = 8'h01;
      17'd38371: data = 8'h04;
      17'd38372: data = 8'h00;
      17'd38373: data = 8'hfa;
      17'd38374: data = 8'hf1;
      17'd38375: data = 8'hf5;
      17'd38376: data = 8'hfe;
      17'd38377: data = 8'hfc;
      17'd38378: data = 8'hf4;
      17'd38379: data = 8'hef;
      17'd38380: data = 8'hf4;
      17'd38381: data = 8'hfa;
      17'd38382: data = 8'hfd;
      17'd38383: data = 8'hfc;
      17'd38384: data = 8'hf4;
      17'd38385: data = 8'hed;
      17'd38386: data = 8'hef;
      17'd38387: data = 8'hf5;
      17'd38388: data = 8'hfc;
      17'd38389: data = 8'hfd;
      17'd38390: data = 8'hf5;
      17'd38391: data = 8'hf4;
      17'd38392: data = 8'hfc;
      17'd38393: data = 8'hf9;
      17'd38394: data = 8'hf2;
      17'd38395: data = 8'hf6;
      17'd38396: data = 8'hf5;
      17'd38397: data = 8'hf1;
      17'd38398: data = 8'hf9;
      17'd38399: data = 8'hf9;
      17'd38400: data = 8'hef;
      17'd38401: data = 8'hfe;
      17'd38402: data = 8'h04;
      17'd38403: data = 8'hf5;
      17'd38404: data = 8'hf2;
      17'd38405: data = 8'hf9;
      17'd38406: data = 8'hfe;
      17'd38407: data = 8'h04;
      17'd38408: data = 8'h04;
      17'd38409: data = 8'h04;
      17'd38410: data = 8'hfd;
      17'd38411: data = 8'hf5;
      17'd38412: data = 8'h00;
      17'd38413: data = 8'h01;
      17'd38414: data = 8'h09;
      17'd38415: data = 8'h11;
      17'd38416: data = 8'hfd;
      17'd38417: data = 8'hf1;
      17'd38418: data = 8'hfe;
      17'd38419: data = 8'h0c;
      17'd38420: data = 8'h11;
      17'd38421: data = 8'h0c;
      17'd38422: data = 8'h01;
      17'd38423: data = 8'hf6;
      17'd38424: data = 8'hf5;
      17'd38425: data = 8'h0a;
      17'd38426: data = 8'h1a;
      17'd38427: data = 8'h11;
      17'd38428: data = 8'hf5;
      17'd38429: data = 8'heb;
      17'd38430: data = 8'h02;
      17'd38431: data = 8'h12;
      17'd38432: data = 8'h0c;
      17'd38433: data = 8'hfe;
      17'd38434: data = 8'hed;
      17'd38435: data = 8'hf4;
      17'd38436: data = 8'h0c;
      17'd38437: data = 8'h13;
      17'd38438: data = 8'hf6;
      17'd38439: data = 8'heb;
      17'd38440: data = 8'h02;
      17'd38441: data = 8'h05;
      17'd38442: data = 8'hfa;
      17'd38443: data = 8'h02;
      17'd38444: data = 8'hfd;
      17'd38445: data = 8'hf9;
      17'd38446: data = 8'h06;
      17'd38447: data = 8'hf9;
      17'd38448: data = 8'hf9;
      17'd38449: data = 8'h09;
      17'd38450: data = 8'h02;
      17'd38451: data = 8'h01;
      17'd38452: data = 8'hfc;
      17'd38453: data = 8'hf4;
      17'd38454: data = 8'h02;
      17'd38455: data = 8'h06;
      17'd38456: data = 8'h05;
      17'd38457: data = 8'hf5;
      17'd38458: data = 8'he5;
      17'd38459: data = 8'h01;
      17'd38460: data = 8'h09;
      17'd38461: data = 8'hf6;
      17'd38462: data = 8'hfe;
      17'd38463: data = 8'h05;
      17'd38464: data = 8'hf5;
      17'd38465: data = 8'hf9;
      17'd38466: data = 8'h0c;
      17'd38467: data = 8'h00;
      17'd38468: data = 8'hfe;
      17'd38469: data = 8'h0a;
      17'd38470: data = 8'hfa;
      17'd38471: data = 8'hfd;
      17'd38472: data = 8'h1a;
      17'd38473: data = 8'h02;
      17'd38474: data = 8'heb;
      17'd38475: data = 8'hfd;
      17'd38476: data = 8'h0a;
      17'd38477: data = 8'h0d;
      17'd38478: data = 8'h05;
      17'd38479: data = 8'h01;
      17'd38480: data = 8'hf2;
      17'd38481: data = 8'hfc;
      17'd38482: data = 8'h0e;
      17'd38483: data = 8'h0a;
      17'd38484: data = 8'hfe;
      17'd38485: data = 8'hfc;
      17'd38486: data = 8'hf4;
      17'd38487: data = 8'hfe;
      17'd38488: data = 8'h26;
      17'd38489: data = 8'h04;
      17'd38490: data = 8'hc6;
      17'd38491: data = 8'h00;
      17'd38492: data = 8'h29;
      17'd38493: data = 8'h01;
      17'd38494: data = 8'hfe;
      17'd38495: data = 8'hdb;
      17'd38496: data = 8'hca;
      17'd38497: data = 8'h3a;
      17'd38498: data = 8'h1c;
      17'd38499: data = 8'hdc;
      17'd38500: data = 8'h04;
      17'd38501: data = 8'hcb;
      17'd38502: data = 8'hfd;
      17'd38503: data = 8'h47;
      17'd38504: data = 8'heb;
      17'd38505: data = 8'he4;
      17'd38506: data = 8'h12;
      17'd38507: data = 8'hfc;
      17'd38508: data = 8'h0e;
      17'd38509: data = 8'h0a;
      17'd38510: data = 8'hf4;
      17'd38511: data = 8'h09;
      17'd38512: data = 8'h22;
      17'd38513: data = 8'h04;
      17'd38514: data = 8'hef;
      17'd38515: data = 8'h19;
      17'd38516: data = 8'h00;
      17'd38517: data = 8'h12;
      17'd38518: data = 8'h23;
      17'd38519: data = 8'hd6;
      17'd38520: data = 8'h0a;
      17'd38521: data = 8'h33;
      17'd38522: data = 8'h0a;
      17'd38523: data = 8'h05;
      17'd38524: data = 8'hed;
      17'd38525: data = 8'hfa;
      17'd38526: data = 8'h27;
      17'd38527: data = 8'h5d;
      17'd38528: data = 8'heb;
      17'd38529: data = 8'haa;
      17'd38530: data = 8'h3c;
      17'd38531: data = 8'h1a;
      17'd38532: data = 8'h00;
      17'd38533: data = 8'h3c;
      17'd38534: data = 8'he3;
      17'd38535: data = 8'hc6;
      17'd38536: data = 8'h3c;
      17'd38537: data = 8'h27;
      17'd38538: data = 8'hdc;
      17'd38539: data = 8'h01;
      17'd38540: data = 8'h15;
      17'd38541: data = 8'h13;
      17'd38542: data = 8'h0c;
      17'd38543: data = 8'hef;
      17'd38544: data = 8'h05;
      17'd38545: data = 8'h1f;
      17'd38546: data = 8'h02;
      17'd38547: data = 8'h0c;
      17'd38548: data = 8'h01;
      17'd38549: data = 8'hfc;
      17'd38550: data = 8'h1a;
      17'd38551: data = 8'h00;
      17'd38552: data = 8'hf9;
      17'd38553: data = 8'h09;
      17'd38554: data = 8'h00;
      17'd38555: data = 8'h12;
      17'd38556: data = 8'h24;
      17'd38557: data = 8'hd8;
      17'd38558: data = 8'hde;
      17'd38559: data = 8'h19;
      17'd38560: data = 8'h1e;
      17'd38561: data = 8'h35;
      17'd38562: data = 8'hd1;
      17'd38563: data = 8'hb8;
      17'd38564: data = 8'h29;
      17'd38565: data = 8'h29;
      17'd38566: data = 8'h22;
      17'd38567: data = 8'hed;
      17'd38568: data = 8'ha2;
      17'd38569: data = 8'h0d;
      17'd38570: data = 8'h56;
      17'd38571: data = 8'h12;
      17'd38572: data = 8'hdb;
      17'd38573: data = 8'hc6;
      17'd38574: data = 8'hfc;
      17'd38575: data = 8'h35;
      17'd38576: data = 8'h2f;
      17'd38577: data = 8'he7;
      17'd38578: data = 8'hd6;
      17'd38579: data = 8'he9;
      17'd38580: data = 8'h22;
      17'd38581: data = 8'h43;
      17'd38582: data = 8'hda;
      17'd38583: data = 8'hda;
      17'd38584: data = 8'h0d;
      17'd38585: data = 8'h02;
      17'd38586: data = 8'h2b;
      17'd38587: data = 8'h01;
      17'd38588: data = 8'hb9;
      17'd38589: data = 8'h12;
      17'd38590: data = 8'h1e;
      17'd38591: data = 8'hfa;
      17'd38592: data = 8'h00;
      17'd38593: data = 8'he0;
      17'd38594: data = 8'hfa;
      17'd38595: data = 8'h11;
      17'd38596: data = 8'h13;
      17'd38597: data = 8'he0;
      17'd38598: data = 8'hcb;
      17'd38599: data = 8'h23;
      17'd38600: data = 8'h34;
      17'd38601: data = 8'hc4;
      17'd38602: data = 8'hd5;
      17'd38603: data = 8'h13;
      17'd38604: data = 8'hf6;
      17'd38605: data = 8'h22;
      17'd38606: data = 8'h02;
      17'd38607: data = 8'hab;
      17'd38608: data = 8'h00;
      17'd38609: data = 8'h31;
      17'd38610: data = 8'he2;
      17'd38611: data = 8'hf6;
      17'd38612: data = 8'h00;
      17'd38613: data = 8'he0;
      17'd38614: data = 8'h02;
      17'd38615: data = 8'h0d;
      17'd38616: data = 8'hef;
      17'd38617: data = 8'h01;
      17'd38618: data = 8'he9;
      17'd38619: data = 8'hf1;
      17'd38620: data = 8'h1b;
      17'd38621: data = 8'he4;
      17'd38622: data = 8'hfa;
      17'd38623: data = 8'h06;
      17'd38624: data = 8'he0;
      17'd38625: data = 8'h09;
      17'd38626: data = 8'hfd;
      17'd38627: data = 8'hef;
      17'd38628: data = 8'h0d;
      17'd38629: data = 8'h02;
      17'd38630: data = 8'hd1;
      17'd38631: data = 8'hfc;
      17'd38632: data = 8'h24;
      17'd38633: data = 8'hec;
      17'd38634: data = 8'hf5;
      17'd38635: data = 8'hf4;
      17'd38636: data = 8'he3;
      17'd38637: data = 8'h02;
      17'd38638: data = 8'h16;
      17'd38639: data = 8'hf4;
      17'd38640: data = 8'hd5;
      17'd38641: data = 8'hef;
      17'd38642: data = 8'h13;
      17'd38643: data = 8'h13;
      17'd38644: data = 8'he3;
      17'd38645: data = 8'hd3;
      17'd38646: data = 8'hfd;
      17'd38647: data = 8'h15;
      17'd38648: data = 8'h12;
      17'd38649: data = 8'he2;
      17'd38650: data = 8'hd8;
      17'd38651: data = 8'h02;
      17'd38652: data = 8'h06;
      17'd38653: data = 8'h0d;
      17'd38654: data = 8'hec;
      17'd38655: data = 8'he9;
      17'd38656: data = 8'h0a;
      17'd38657: data = 8'hf6;
      17'd38658: data = 8'hfd;
      17'd38659: data = 8'h05;
      17'd38660: data = 8'hf2;
      17'd38661: data = 8'hf5;
      17'd38662: data = 8'hf9;
      17'd38663: data = 8'hfd;
      17'd38664: data = 8'hfd;
      17'd38665: data = 8'hf6;
      17'd38666: data = 8'h05;
      17'd38667: data = 8'hef;
      17'd38668: data = 8'heb;
      17'd38669: data = 8'h06;
      17'd38670: data = 8'hf1;
      17'd38671: data = 8'h01;
      17'd38672: data = 8'h15;
      17'd38673: data = 8'hde;
      17'd38674: data = 8'hd8;
      17'd38675: data = 8'h0a;
      17'd38676: data = 8'h12;
      17'd38677: data = 8'h0d;
      17'd38678: data = 8'hf9;
      17'd38679: data = 8'hc5;
      17'd38680: data = 8'hf1;
      17'd38681: data = 8'h24;
      17'd38682: data = 8'h01;
      17'd38683: data = 8'hec;
      17'd38684: data = 8'hf4;
      17'd38685: data = 8'he7;
      17'd38686: data = 8'h0e;
      17'd38687: data = 8'h0e;
      17'd38688: data = 8'hd8;
      17'd38689: data = 8'h0d;
      17'd38690: data = 8'h09;
      17'd38691: data = 8'hda;
      17'd38692: data = 8'h06;
      17'd38693: data = 8'h12;
      17'd38694: data = 8'hf1;
      17'd38695: data = 8'hf2;
      17'd38696: data = 8'hfd;
      17'd38697: data = 8'hfa;
      17'd38698: data = 8'hfd;
      17'd38699: data = 8'hfc;
      17'd38700: data = 8'hec;
      17'd38701: data = 8'hf9;
      17'd38702: data = 8'hfe;
      17'd38703: data = 8'hf4;
      17'd38704: data = 8'h01;
      17'd38705: data = 8'h02;
      17'd38706: data = 8'hf9;
      17'd38707: data = 8'hf4;
      17'd38708: data = 8'hf9;
      17'd38709: data = 8'h0c;
      17'd38710: data = 8'h00;
      17'd38711: data = 8'hf6;
      17'd38712: data = 8'h04;
      17'd38713: data = 8'hfc;
      17'd38714: data = 8'hfe;
      17'd38715: data = 8'h05;
      17'd38716: data = 8'hfe;
      17'd38717: data = 8'h06;
      17'd38718: data = 8'hf9;
      17'd38719: data = 8'hfd;
      17'd38720: data = 8'h11;
      17'd38721: data = 8'h04;
      17'd38722: data = 8'hfc;
      17'd38723: data = 8'h0c;
      17'd38724: data = 8'hfd;
      17'd38725: data = 8'hfa;
      17'd38726: data = 8'h15;
      17'd38727: data = 8'hfd;
      17'd38728: data = 8'hfa;
      17'd38729: data = 8'h04;
      17'd38730: data = 8'hfc;
      17'd38731: data = 8'h0e;
      17'd38732: data = 8'h04;
      17'd38733: data = 8'hfc;
      17'd38734: data = 8'hfd;
      17'd38735: data = 8'hf2;
      17'd38736: data = 8'h05;
      17'd38737: data = 8'h26;
      17'd38738: data = 8'hf6;
      17'd38739: data = 8'he5;
      17'd38740: data = 8'h12;
      17'd38741: data = 8'h02;
      17'd38742: data = 8'h01;
      17'd38743: data = 8'h0a;
      17'd38744: data = 8'h06;
      17'd38745: data = 8'h05;
      17'd38746: data = 8'hef;
      17'd38747: data = 8'hfd;
      17'd38748: data = 8'h15;
      17'd38749: data = 8'h01;
      17'd38750: data = 8'h0c;
      17'd38751: data = 8'h05;
      17'd38752: data = 8'he9;
      17'd38753: data = 8'h04;
      17'd38754: data = 8'h16;
      17'd38755: data = 8'h0d;
      17'd38756: data = 8'hf5;
      17'd38757: data = 8'hfc;
      17'd38758: data = 8'h02;
      17'd38759: data = 8'hfe;
      17'd38760: data = 8'h1f;
      17'd38761: data = 8'h0a;
      17'd38762: data = 8'hf1;
      17'd38763: data = 8'hfa;
      17'd38764: data = 8'hfa;
      17'd38765: data = 8'h1a;
      17'd38766: data = 8'h1b;
      17'd38767: data = 8'hef;
      17'd38768: data = 8'hef;
      17'd38769: data = 8'h01;
      17'd38770: data = 8'h0d;
      17'd38771: data = 8'h22;
      17'd38772: data = 8'hfc;
      17'd38773: data = 8'he7;
      17'd38774: data = 8'h0e;
      17'd38775: data = 8'h05;
      17'd38776: data = 8'h0a;
      17'd38777: data = 8'h1a;
      17'd38778: data = 8'h02;
      17'd38779: data = 8'hfa;
      17'd38780: data = 8'hfc;
      17'd38781: data = 8'h16;
      17'd38782: data = 8'h1f;
      17'd38783: data = 8'h00;
      17'd38784: data = 8'hef;
      17'd38785: data = 8'h00;
      17'd38786: data = 8'h23;
      17'd38787: data = 8'h0a;
      17'd38788: data = 8'hfc;
      17'd38789: data = 8'h05;
      17'd38790: data = 8'hed;
      17'd38791: data = 8'h02;
      17'd38792: data = 8'h35;
      17'd38793: data = 8'h0c;
      17'd38794: data = 8'hc9;
      17'd38795: data = 8'hf5;
      17'd38796: data = 8'h1f;
      17'd38797: data = 8'h15;
      17'd38798: data = 8'h1b;
      17'd38799: data = 8'he3;
      17'd38800: data = 8'hc6;
      17'd38801: data = 8'h24;
      17'd38802: data = 8'h26;
      17'd38803: data = 8'hf9;
      17'd38804: data = 8'hfa;
      17'd38805: data = 8'hdb;
      17'd38806: data = 8'hfe;
      17'd38807: data = 8'h2c;
      17'd38808: data = 8'h0c;
      17'd38809: data = 8'he4;
      17'd38810: data = 8'he7;
      17'd38811: data = 8'h1e;
      17'd38812: data = 8'h0c;
      17'd38813: data = 8'hf4;
      17'd38814: data = 8'h09;
      17'd38815: data = 8'hfe;
      17'd38816: data = 8'hf6;
      17'd38817: data = 8'h1a;
      17'd38818: data = 8'h1c;
      17'd38819: data = 8'hd8;
      17'd38820: data = 8'hed;
      17'd38821: data = 8'h2b;
      17'd38822: data = 8'h0e;
      17'd38823: data = 8'hf4;
      17'd38824: data = 8'hf1;
      17'd38825: data = 8'h02;
      17'd38826: data = 8'h0a;
      17'd38827: data = 8'hf6;
      17'd38828: data = 8'h0e;
      17'd38829: data = 8'h00;
      17'd38830: data = 8'he7;
      17'd38831: data = 8'h0a;
      17'd38832: data = 8'h04;
      17'd38833: data = 8'h02;
      17'd38834: data = 8'hfe;
      17'd38835: data = 8'h05;
      17'd38836: data = 8'h00;
      17'd38837: data = 8'he3;
      17'd38838: data = 8'h05;
      17'd38839: data = 8'h0c;
      17'd38840: data = 8'h33;
      17'd38841: data = 8'he2;
      17'd38842: data = 8'hb4;
      17'd38843: data = 8'h33;
      17'd38844: data = 8'h2d;
      17'd38845: data = 8'hec;
      17'd38846: data = 8'hed;
      17'd38847: data = 8'hf6;
      17'd38848: data = 8'hfc;
      17'd38849: data = 8'h29;
      17'd38850: data = 8'h01;
      17'd38851: data = 8'he9;
      17'd38852: data = 8'h04;
      17'd38853: data = 8'hfd;
      17'd38854: data = 8'h01;
      17'd38855: data = 8'h0c;
      17'd38856: data = 8'hfe;
      17'd38857: data = 8'hf9;
      17'd38858: data = 8'hf1;
      17'd38859: data = 8'hfc;
      17'd38860: data = 8'h16;
      17'd38861: data = 8'h00;
      17'd38862: data = 8'hec;
      17'd38863: data = 8'hf2;
      17'd38864: data = 8'h0c;
      17'd38865: data = 8'h01;
      17'd38866: data = 8'hf2;
      17'd38867: data = 8'h09;
      17'd38868: data = 8'hf9;
      17'd38869: data = 8'hfa;
      17'd38870: data = 8'hf5;
      17'd38871: data = 8'h11;
      17'd38872: data = 8'hf5;
      17'd38873: data = 8'he4;
      17'd38874: data = 8'h27;
      17'd38875: data = 8'hf9;
      17'd38876: data = 8'hdb;
      17'd38877: data = 8'h19;
      17'd38878: data = 8'h04;
      17'd38879: data = 8'hef;
      17'd38880: data = 8'h19;
      17'd38881: data = 8'he4;
      17'd38882: data = 8'he3;
      17'd38883: data = 8'h23;
      17'd38884: data = 8'h1b;
      17'd38885: data = 8'he0;
      17'd38886: data = 8'hf1;
      17'd38887: data = 8'h0e;
      17'd38888: data = 8'hfa;
      17'd38889: data = 8'h12;
      17'd38890: data = 8'hf2;
      17'd38891: data = 8'hfa;
      17'd38892: data = 8'h06;
      17'd38893: data = 8'hf6;
      17'd38894: data = 8'h19;
      17'd38895: data = 8'hf1;
      17'd38896: data = 8'heb;
      17'd38897: data = 8'h11;
      17'd38898: data = 8'hf6;
      17'd38899: data = 8'h04;
      17'd38900: data = 8'hfc;
      17'd38901: data = 8'he4;
      17'd38902: data = 8'h0a;
      17'd38903: data = 8'hf6;
      17'd38904: data = 8'h06;
      17'd38905: data = 8'hf9;
      17'd38906: data = 8'he5;
      17'd38907: data = 8'h12;
      17'd38908: data = 8'hf4;
      17'd38909: data = 8'hf2;
      17'd38910: data = 8'hfa;
      17'd38911: data = 8'hfc;
      17'd38912: data = 8'h19;
      17'd38913: data = 8'hf4;
      17'd38914: data = 8'he0;
      17'd38915: data = 8'hf5;
      17'd38916: data = 8'h0d;
      17'd38917: data = 8'h1e;
      17'd38918: data = 8'he4;
      17'd38919: data = 8'hca;
      17'd38920: data = 8'h0d;
      17'd38921: data = 8'h1a;
      17'd38922: data = 8'h0c;
      17'd38923: data = 8'h01;
      17'd38924: data = 8'hc1;
      17'd38925: data = 8'hf4;
      17'd38926: data = 8'h33;
      17'd38927: data = 8'h09;
      17'd38928: data = 8'hf1;
      17'd38929: data = 8'hda;
      17'd38930: data = 8'hf6;
      17'd38931: data = 8'h11;
      17'd38932: data = 8'h13;
      17'd38933: data = 8'hfd;
      17'd38934: data = 8'hda;
      17'd38935: data = 8'hed;
      17'd38936: data = 8'h01;
      17'd38937: data = 8'h23;
      17'd38938: data = 8'hfd;
      17'd38939: data = 8'hc4;
      17'd38940: data = 8'h11;
      17'd38941: data = 8'h11;
      17'd38942: data = 8'hf5;
      17'd38943: data = 8'h0c;
      17'd38944: data = 8'he2;
      17'd38945: data = 8'hfa;
      17'd38946: data = 8'hf9;
      17'd38947: data = 8'h0c;
      17'd38948: data = 8'h0d;
      17'd38949: data = 8'hdb;
      17'd38950: data = 8'h12;
      17'd38951: data = 8'hfc;
      17'd38952: data = 8'he7;
      17'd38953: data = 8'h09;
      17'd38954: data = 8'hf2;
      17'd38955: data = 8'h11;
      17'd38956: data = 8'h0e;
      17'd38957: data = 8'hd5;
      17'd38958: data = 8'hfe;
      17'd38959: data = 8'h19;
      17'd38960: data = 8'h00;
      17'd38961: data = 8'hfe;
      17'd38962: data = 8'he4;
      17'd38963: data = 8'h06;
      17'd38964: data = 8'h23;
      17'd38965: data = 8'hd2;
      17'd38966: data = 8'hf2;
      17'd38967: data = 8'h2f;
      17'd38968: data = 8'he5;
      17'd38969: data = 8'hfa;
      17'd38970: data = 8'h29;
      17'd38971: data = 8'hce;
      17'd38972: data = 8'hec;
      17'd38973: data = 8'h3a;
      17'd38974: data = 8'h04;
      17'd38975: data = 8'hd5;
      17'd38976: data = 8'hf4;
      17'd38977: data = 8'h16;
      17'd38978: data = 8'h04;
      17'd38979: data = 8'h04;
      17'd38980: data = 8'hf6;
      17'd38981: data = 8'he0;
      17'd38982: data = 8'h09;
      17'd38983: data = 8'h23;
      17'd38984: data = 8'hfc;
      17'd38985: data = 8'he9;
      17'd38986: data = 8'h06;
      17'd38987: data = 8'h09;
      17'd38988: data = 8'h06;
      17'd38989: data = 8'hfc;
      17'd38990: data = 8'hf6;
      17'd38991: data = 8'h05;
      17'd38992: data = 8'hfd;
      17'd38993: data = 8'h1a;
      17'd38994: data = 8'he7;
      17'd38995: data = 8'hd8;
      17'd38996: data = 8'h2f;
      17'd38997: data = 8'h22;
      17'd38998: data = 8'hd5;
      17'd38999: data = 8'he4;
      17'd39000: data = 8'h12;
      17'd39001: data = 8'hfc;
      17'd39002: data = 8'h15;
      17'd39003: data = 8'hf6;
      17'd39004: data = 8'hde;
      17'd39005: data = 8'h09;
      17'd39006: data = 8'h05;
      17'd39007: data = 8'hfd;
      17'd39008: data = 8'hf4;
      17'd39009: data = 8'hfd;
      17'd39010: data = 8'h00;
      17'd39011: data = 8'hf4;
      17'd39012: data = 8'h15;
      17'd39013: data = 8'h01;
      17'd39014: data = 8'hf2;
      17'd39015: data = 8'h09;
      17'd39016: data = 8'hec;
      17'd39017: data = 8'h1a;
      17'd39018: data = 8'hfd;
      17'd39019: data = 8'hde;
      17'd39020: data = 8'h1b;
      17'd39021: data = 8'hfa;
      17'd39022: data = 8'hfe;
      17'd39023: data = 8'h09;
      17'd39024: data = 8'hf2;
      17'd39025: data = 8'h05;
      17'd39026: data = 8'h0a;
      17'd39027: data = 8'hf1;
      17'd39028: data = 8'h0e;
      17'd39029: data = 8'h16;
      17'd39030: data = 8'hdc;
      17'd39031: data = 8'hfa;
      17'd39032: data = 8'h19;
      17'd39033: data = 8'h0a;
      17'd39034: data = 8'h0e;
      17'd39035: data = 8'hef;
      17'd39036: data = 8'hf5;
      17'd39037: data = 8'hfc;
      17'd39038: data = 8'h12;
      17'd39039: data = 8'h1c;
      17'd39040: data = 8'he4;
      17'd39041: data = 8'h04;
      17'd39042: data = 8'hf5;
      17'd39043: data = 8'h01;
      17'd39044: data = 8'h27;
      17'd39045: data = 8'hfa;
      17'd39046: data = 8'hed;
      17'd39047: data = 8'hf9;
      17'd39048: data = 8'h16;
      17'd39049: data = 8'h19;
      17'd39050: data = 8'hf2;
      17'd39051: data = 8'h05;
      17'd39052: data = 8'h05;
      17'd39053: data = 8'hf5;
      17'd39054: data = 8'h19;
      17'd39055: data = 8'h06;
      17'd39056: data = 8'heb;
      17'd39057: data = 8'hfa;
      17'd39058: data = 8'h1a;
      17'd39059: data = 8'h04;
      17'd39060: data = 8'he2;
      17'd39061: data = 8'h15;
      17'd39062: data = 8'h12;
      17'd39063: data = 8'hd1;
      17'd39064: data = 8'h13;
      17'd39065: data = 8'h1b;
      17'd39066: data = 8'hd2;
      17'd39067: data = 8'h15;
      17'd39068: data = 8'h00;
      17'd39069: data = 8'hf2;
      17'd39070: data = 8'h0a;
      17'd39071: data = 8'he5;
      17'd39072: data = 8'h12;
      17'd39073: data = 8'h11;
      17'd39074: data = 8'hef;
      17'd39075: data = 8'he7;
      17'd39076: data = 8'h06;
      17'd39077: data = 8'h1f;
      17'd39078: data = 8'hf6;
      17'd39079: data = 8'hf4;
      17'd39080: data = 8'h01;
      17'd39081: data = 8'hfa;
      17'd39082: data = 8'h13;
      17'd39083: data = 8'h0d;
      17'd39084: data = 8'heb;
      17'd39085: data = 8'hf6;
      17'd39086: data = 8'h06;
      17'd39087: data = 8'h1b;
      17'd39088: data = 8'h0c;
      17'd39089: data = 8'he2;
      17'd39090: data = 8'h01;
      17'd39091: data = 8'h09;
      17'd39092: data = 8'hfe;
      17'd39093: data = 8'h1a;
      17'd39094: data = 8'h0c;
      17'd39095: data = 8'hdc;
      17'd39096: data = 8'hf5;
      17'd39097: data = 8'h2b;
      17'd39098: data = 8'h06;
      17'd39099: data = 8'he5;
      17'd39100: data = 8'hfa;
      17'd39101: data = 8'h04;
      17'd39102: data = 8'h09;
      17'd39103: data = 8'h1a;
      17'd39104: data = 8'hed;
      17'd39105: data = 8'he5;
      17'd39106: data = 8'h13;
      17'd39107: data = 8'h11;
      17'd39108: data = 8'h09;
      17'd39109: data = 8'he5;
      17'd39110: data = 8'hfc;
      17'd39111: data = 8'h19;
      17'd39112: data = 8'he9;
      17'd39113: data = 8'h01;
      17'd39114: data = 8'h0d;
      17'd39115: data = 8'heb;
      17'd39116: data = 8'h04;
      17'd39117: data = 8'h00;
      17'd39118: data = 8'h00;
      17'd39119: data = 8'h00;
      17'd39120: data = 8'hf6;
      17'd39121: data = 8'h04;
      17'd39122: data = 8'h05;
      17'd39123: data = 8'h09;
      17'd39124: data = 8'hf4;
      17'd39125: data = 8'hf9;
      17'd39126: data = 8'h0d;
      17'd39127: data = 8'hfc;
      17'd39128: data = 8'hf4;
      17'd39129: data = 8'h22;
      17'd39130: data = 8'hf1;
      17'd39131: data = 8'hec;
      17'd39132: data = 8'h26;
      17'd39133: data = 8'heb;
      17'd39134: data = 8'hf9;
      17'd39135: data = 8'h11;
      17'd39136: data = 8'hec;
      17'd39137: data = 8'h1a;
      17'd39138: data = 8'h01;
      17'd39139: data = 8'hd8;
      17'd39140: data = 8'h12;
      17'd39141: data = 8'h15;
      17'd39142: data = 8'he3;
      17'd39143: data = 8'hf9;
      17'd39144: data = 8'h22;
      17'd39145: data = 8'hf1;
      17'd39146: data = 8'hf4;
      17'd39147: data = 8'h0c;
      17'd39148: data = 8'he9;
      17'd39149: data = 8'h11;
      17'd39150: data = 8'h13;
      17'd39151: data = 8'hec;
      17'd39152: data = 8'hfe;
      17'd39153: data = 8'h00;
      17'd39154: data = 8'hf6;
      17'd39155: data = 8'h13;
      17'd39156: data = 8'hfe;
      17'd39157: data = 8'he4;
      17'd39158: data = 8'h11;
      17'd39159: data = 8'h09;
      17'd39160: data = 8'heb;
      17'd39161: data = 8'hf2;
      17'd39162: data = 8'h0e;
      17'd39163: data = 8'hed;
      17'd39164: data = 8'hf5;
      17'd39165: data = 8'h1e;
      17'd39166: data = 8'he7;
      17'd39167: data = 8'he9;
      17'd39168: data = 8'h05;
      17'd39169: data = 8'hfe;
      17'd39170: data = 8'h02;
      17'd39171: data = 8'hfc;
      17'd39172: data = 8'hf1;
      17'd39173: data = 8'hf9;
      17'd39174: data = 8'hfc;
      17'd39175: data = 8'h0c;
      17'd39176: data = 8'hfc;
      17'd39177: data = 8'hec;
      17'd39178: data = 8'h0c;
      17'd39179: data = 8'hfc;
      17'd39180: data = 8'hf2;
      17'd39181: data = 8'h0c;
      17'd39182: data = 8'he9;
      17'd39183: data = 8'h0a;
      17'd39184: data = 8'h1b;
      17'd39185: data = 8'hec;
      17'd39186: data = 8'hef;
      17'd39187: data = 8'h02;
      17'd39188: data = 8'hfe;
      17'd39189: data = 8'h0e;
      17'd39190: data = 8'h19;
      17'd39191: data = 8'he4;
      17'd39192: data = 8'hf1;
      17'd39193: data = 8'h0d;
      17'd39194: data = 8'h0e;
      17'd39195: data = 8'h06;
      17'd39196: data = 8'hf5;
      17'd39197: data = 8'hfd;
      17'd39198: data = 8'h05;
      17'd39199: data = 8'h05;
      17'd39200: data = 8'hf5;
      17'd39201: data = 8'hfc;
      17'd39202: data = 8'h0e;
      17'd39203: data = 8'hf4;
      17'd39204: data = 8'h00;
      17'd39205: data = 8'h09;
      17'd39206: data = 8'he5;
      17'd39207: data = 8'h02;
      17'd39208: data = 8'h11;
      17'd39209: data = 8'hfc;
      17'd39210: data = 8'hf9;
      17'd39211: data = 8'hf5;
      17'd39212: data = 8'hf9;
      17'd39213: data = 8'h13;
      17'd39214: data = 8'h13;
      17'd39215: data = 8'hd6;
      17'd39216: data = 8'hf9;
      17'd39217: data = 8'h15;
      17'd39218: data = 8'hed;
      17'd39219: data = 8'h0a;
      17'd39220: data = 8'hfc;
      17'd39221: data = 8'he2;
      17'd39222: data = 8'h13;
      17'd39223: data = 8'h06;
      17'd39224: data = 8'hef;
      17'd39225: data = 8'h04;
      17'd39226: data = 8'hf2;
      17'd39227: data = 8'hf4;
      17'd39228: data = 8'h26;
      17'd39229: data = 8'h02;
      17'd39230: data = 8'hd5;
      17'd39231: data = 8'h0c;
      17'd39232: data = 8'h11;
      17'd39233: data = 8'hfa;
      17'd39234: data = 8'h0e;
      17'd39235: data = 8'hef;
      17'd39236: data = 8'hd8;
      17'd39237: data = 8'h2b;
      17'd39238: data = 8'h0d;
      17'd39239: data = 8'hda;
      17'd39240: data = 8'h15;
      17'd39241: data = 8'he9;
      17'd39242: data = 8'hf4;
      17'd39243: data = 8'h3a;
      17'd39244: data = 8'hf2;
      17'd39245: data = 8'hd2;
      17'd39246: data = 8'h15;
      17'd39247: data = 8'h04;
      17'd39248: data = 8'h11;
      17'd39249: data = 8'h11;
      17'd39250: data = 8'hda;
      17'd39251: data = 8'hf9;
      17'd39252: data = 8'h1e;
      17'd39253: data = 8'h0a;
      17'd39254: data = 8'he7;
      17'd39255: data = 8'hfa;
      17'd39256: data = 8'h00;
      17'd39257: data = 8'h12;
      17'd39258: data = 8'h06;
      17'd39259: data = 8'he3;
      17'd39260: data = 8'hfa;
      17'd39261: data = 8'h06;
      17'd39262: data = 8'h06;
      17'd39263: data = 8'h04;
      17'd39264: data = 8'he0;
      17'd39265: data = 8'hef;
      17'd39266: data = 8'h1c;
      17'd39267: data = 8'hfc;
      17'd39268: data = 8'hed;
      17'd39269: data = 8'h06;
      17'd39270: data = 8'he5;
      17'd39271: data = 8'hfd;
      17'd39272: data = 8'h1f;
      17'd39273: data = 8'he0;
      17'd39274: data = 8'hfd;
      17'd39275: data = 8'hf9;
      17'd39276: data = 8'hfa;
      17'd39277: data = 8'h1e;
      17'd39278: data = 8'he2;
      17'd39279: data = 8'hf1;
      17'd39280: data = 8'h06;
      17'd39281: data = 8'h01;
      17'd39282: data = 8'h0d;
      17'd39283: data = 8'he0;
      17'd39284: data = 8'hfc;
      17'd39285: data = 8'h1b;
      17'd39286: data = 8'hf2;
      17'd39287: data = 8'h01;
      17'd39288: data = 8'h01;
      17'd39289: data = 8'hf9;
      17'd39290: data = 8'h06;
      17'd39291: data = 8'h0c;
      17'd39292: data = 8'h00;
      17'd39293: data = 8'hf9;
      17'd39294: data = 8'h00;
      17'd39295: data = 8'hfc;
      17'd39296: data = 8'h16;
      17'd39297: data = 8'h15;
      17'd39298: data = 8'hd2;
      17'd39299: data = 8'h04;
      17'd39300: data = 8'h1a;
      17'd39301: data = 8'he4;
      17'd39302: data = 8'h11;
      17'd39303: data = 8'h0c;
      17'd39304: data = 8'heb;
      17'd39305: data = 8'hf5;
      17'd39306: data = 8'h16;
      17'd39307: data = 8'h0d;
      17'd39308: data = 8'he4;
      17'd39309: data = 8'h00;
      17'd39310: data = 8'h0a;
      17'd39311: data = 8'h00;
      17'd39312: data = 8'h04;
      17'd39313: data = 8'heb;
      17'd39314: data = 8'hf9;
      17'd39315: data = 8'h23;
      17'd39316: data = 8'h02;
      17'd39317: data = 8'hd8;
      17'd39318: data = 8'hfc;
      17'd39319: data = 8'h0e;
      17'd39320: data = 8'h09;
      17'd39321: data = 8'hfd;
      17'd39322: data = 8'he5;
      17'd39323: data = 8'hfc;
      17'd39324: data = 8'h0c;
      17'd39325: data = 8'h1c;
      17'd39326: data = 8'hf4;
      17'd39327: data = 8'he0;
      17'd39328: data = 8'h06;
      17'd39329: data = 8'h01;
      17'd39330: data = 8'h0e;
      17'd39331: data = 8'h0c;
      17'd39332: data = 8'he7;
      17'd39333: data = 8'hfd;
      17'd39334: data = 8'hf6;
      17'd39335: data = 8'h26;
      17'd39336: data = 8'h16;
      17'd39337: data = 8'hb4;
      17'd39338: data = 8'h09;
      17'd39339: data = 8'h22;
      17'd39340: data = 8'h02;
      17'd39341: data = 8'h09;
      17'd39342: data = 8'hdb;
      17'd39343: data = 8'hef;
      17'd39344: data = 8'h22;
      17'd39345: data = 8'h13;
      17'd39346: data = 8'hf1;
      17'd39347: data = 8'hdb;
      17'd39348: data = 8'h11;
      17'd39349: data = 8'h26;
      17'd39350: data = 8'he3;
      17'd39351: data = 8'h02;
      17'd39352: data = 8'h04;
      17'd39353: data = 8'hf2;
      17'd39354: data = 8'h27;
      17'd39355: data = 8'hfa;
      17'd39356: data = 8'hdc;
      17'd39357: data = 8'h12;
      17'd39358: data = 8'h0d;
      17'd39359: data = 8'hfc;
      17'd39360: data = 8'hfc;
      17'd39361: data = 8'hfc;
      17'd39362: data = 8'h01;
      17'd39363: data = 8'h11;
      17'd39364: data = 8'h09;
      17'd39365: data = 8'he0;
      17'd39366: data = 8'hf5;
      17'd39367: data = 8'h1e;
      17'd39368: data = 8'h0a;
      17'd39369: data = 8'hf1;
      17'd39370: data = 8'hf4;
      17'd39371: data = 8'hf6;
      17'd39372: data = 8'h05;
      17'd39373: data = 8'h19;
      17'd39374: data = 8'hec;
      17'd39375: data = 8'he5;
      17'd39376: data = 8'h0c;
      17'd39377: data = 8'h06;
      17'd39378: data = 8'h02;
      17'd39379: data = 8'hfd;
      17'd39380: data = 8'he4;
      17'd39381: data = 8'h04;
      17'd39382: data = 8'h22;
      17'd39383: data = 8'hfe;
      17'd39384: data = 8'hf1;
      17'd39385: data = 8'he5;
      17'd39386: data = 8'hf5;
      17'd39387: data = 8'h39;
      17'd39388: data = 8'h1a;
      17'd39389: data = 8'hca;
      17'd39390: data = 8'he4;
      17'd39391: data = 8'h12;
      17'd39392: data = 8'h2b;
      17'd39393: data = 8'h0a;
      17'd39394: data = 8'hdc;
      17'd39395: data = 8'he9;
      17'd39396: data = 8'h04;
      17'd39397: data = 8'h22;
      17'd39398: data = 8'h12;
      17'd39399: data = 8'hd6;
      17'd39400: data = 8'hec;
      17'd39401: data = 8'h1c;
      17'd39402: data = 8'h13;
      17'd39403: data = 8'hf5;
      17'd39404: data = 8'he9;
      17'd39405: data = 8'h04;
      17'd39406: data = 8'h0a;
      17'd39407: data = 8'hfd;
      17'd39408: data = 8'h01;
      17'd39409: data = 8'h0a;
      17'd39410: data = 8'hec;
      17'd39411: data = 8'hec;
      17'd39412: data = 8'h13;
      17'd39413: data = 8'h15;
      17'd39414: data = 8'h05;
      17'd39415: data = 8'hd3;
      17'd39416: data = 8'hf6;
      17'd39417: data = 8'h29;
      17'd39418: data = 8'hfc;
      17'd39419: data = 8'hed;
      17'd39420: data = 8'h01;
      17'd39421: data = 8'hf9;
      17'd39422: data = 8'h00;
      17'd39423: data = 8'h0c;
      17'd39424: data = 8'hf2;
      17'd39425: data = 8'h0d;
      17'd39426: data = 8'hf2;
      17'd39427: data = 8'hef;
      17'd39428: data = 8'h12;
      17'd39429: data = 8'hfd;
      17'd39430: data = 8'h0a;
      17'd39431: data = 8'hec;
      17'd39432: data = 8'hfd;
      17'd39433: data = 8'h0e;
      17'd39434: data = 8'hed;
      17'd39435: data = 8'h0a;
      17'd39436: data = 8'h0c;
      17'd39437: data = 8'hd8;
      17'd39438: data = 8'h02;
      17'd39439: data = 8'h1b;
      17'd39440: data = 8'hfd;
      17'd39441: data = 8'hf9;
      17'd39442: data = 8'hf4;
      17'd39443: data = 8'h09;
      17'd39444: data = 8'hfc;
      17'd39445: data = 8'h13;
      17'd39446: data = 8'h05;
      17'd39447: data = 8'he5;
      17'd39448: data = 8'h0c;
      17'd39449: data = 8'h02;
      17'd39450: data = 8'h04;
      17'd39451: data = 8'hf4;
      17'd39452: data = 8'h04;
      17'd39453: data = 8'h1f;
      17'd39454: data = 8'he3;
      17'd39455: data = 8'hed;
      17'd39456: data = 8'h19;
      17'd39457: data = 8'h12;
      17'd39458: data = 8'h01;
      17'd39459: data = 8'hed;
      17'd39460: data = 8'hf9;
      17'd39461: data = 8'h0a;
      17'd39462: data = 8'h00;
      17'd39463: data = 8'h19;
      17'd39464: data = 8'hfd;
      17'd39465: data = 8'hd3;
      17'd39466: data = 8'h19;
      17'd39467: data = 8'h1b;
      17'd39468: data = 8'hf5;
      17'd39469: data = 8'hfe;
      17'd39470: data = 8'hf5;
      17'd39471: data = 8'hed;
      17'd39472: data = 8'h12;
      17'd39473: data = 8'h16;
      17'd39474: data = 8'hec;
      17'd39475: data = 8'hf1;
      17'd39476: data = 8'hf5;
      17'd39477: data = 8'h00;
      17'd39478: data = 8'h1a;
      17'd39479: data = 8'h01;
      17'd39480: data = 8'he2;
      17'd39481: data = 8'hfd;
      17'd39482: data = 8'h0e;
      17'd39483: data = 8'h00;
      17'd39484: data = 8'h00;
      17'd39485: data = 8'h0e;
      17'd39486: data = 8'hf9;
      17'd39487: data = 8'he3;
      17'd39488: data = 8'h12;
      17'd39489: data = 8'h12;
      17'd39490: data = 8'hf1;
      17'd39491: data = 8'hf6;
      17'd39492: data = 8'hfc;
      17'd39493: data = 8'hfd;
      17'd39494: data = 8'h13;
      17'd39495: data = 8'h01;
      17'd39496: data = 8'hf5;
      17'd39497: data = 8'hfa;
      17'd39498: data = 8'hf6;
      17'd39499: data = 8'h0c;
      17'd39500: data = 8'h0d;
      17'd39501: data = 8'hf5;
      17'd39502: data = 8'hed;
      17'd39503: data = 8'h02;
      17'd39504: data = 8'h04;
      17'd39505: data = 8'h02;
      17'd39506: data = 8'hfe;
      17'd39507: data = 8'hfe;
      17'd39508: data = 8'hf9;
      17'd39509: data = 8'h02;
      17'd39510: data = 8'h02;
      17'd39511: data = 8'hfe;
      17'd39512: data = 8'h06;
      17'd39513: data = 8'hf4;
      17'd39514: data = 8'h06;
      17'd39515: data = 8'h01;
      17'd39516: data = 8'hf1;
      17'd39517: data = 8'h06;
      17'd39518: data = 8'h01;
      17'd39519: data = 8'hfc;
      17'd39520: data = 8'h04;
      17'd39521: data = 8'h02;
      17'd39522: data = 8'hf5;
      17'd39523: data = 8'h01;
      17'd39524: data = 8'h04;
      17'd39525: data = 8'heb;
      17'd39526: data = 8'h0c;
      17'd39527: data = 8'h06;
      17'd39528: data = 8'he9;
      17'd39529: data = 8'h09;
      17'd39530: data = 8'hfa;
      17'd39531: data = 8'he9;
      17'd39532: data = 8'h0d;
      17'd39533: data = 8'h15;
      17'd39534: data = 8'hed;
      17'd39535: data = 8'hf1;
      17'd39536: data = 8'h01;
      17'd39537: data = 8'hfd;
      17'd39538: data = 8'h0a;
      17'd39539: data = 8'h05;
      17'd39540: data = 8'hf2;
      17'd39541: data = 8'hf9;
      17'd39542: data = 8'h13;
      17'd39543: data = 8'h00;
      17'd39544: data = 8'hf5;
      17'd39545: data = 8'h01;
      17'd39546: data = 8'h06;
      17'd39547: data = 8'hf9;
      17'd39548: data = 8'h00;
      17'd39549: data = 8'h13;
      17'd39550: data = 8'he4;
      17'd39551: data = 8'h01;
      17'd39552: data = 8'h0d;
      17'd39553: data = 8'hf5;
      17'd39554: data = 8'hfe;
      17'd39555: data = 8'hf4;
      17'd39556: data = 8'h02;
      17'd39557: data = 8'h06;
      17'd39558: data = 8'hf1;
      17'd39559: data = 8'hf9;
      17'd39560: data = 8'h02;
      17'd39561: data = 8'hfe;
      17'd39562: data = 8'h1a;
      17'd39563: data = 8'hec;
      17'd39564: data = 8'he3;
      17'd39565: data = 8'h1a;
      17'd39566: data = 8'h02;
      17'd39567: data = 8'hfc;
      17'd39568: data = 8'h0c;
      17'd39569: data = 8'hf5;
      17'd39570: data = 8'hec;
      17'd39571: data = 8'h0e;
      17'd39572: data = 8'h04;
      17'd39573: data = 8'hfa;
      17'd39574: data = 8'h02;
      17'd39575: data = 8'hef;
      17'd39576: data = 8'hf6;
      17'd39577: data = 8'h19;
      17'd39578: data = 8'hf4;
      17'd39579: data = 8'hf5;
      17'd39580: data = 8'h02;
      17'd39581: data = 8'hfa;
      17'd39582: data = 8'h0c;
      17'd39583: data = 8'he9;
      17'd39584: data = 8'hf5;
      17'd39585: data = 8'h12;
      17'd39586: data = 8'hf5;
      17'd39587: data = 8'hfe;
      17'd39588: data = 8'h06;
      17'd39589: data = 8'he7;
      17'd39590: data = 8'h01;
      17'd39591: data = 8'h12;
      17'd39592: data = 8'hef;
      17'd39593: data = 8'h05;
      17'd39594: data = 8'h0a;
      17'd39595: data = 8'he7;
      17'd39596: data = 8'h01;
      17'd39597: data = 8'h1a;
      17'd39598: data = 8'hfc;
      17'd39599: data = 8'hed;
      17'd39600: data = 8'hfa;
      17'd39601: data = 8'hfa;
      17'd39602: data = 8'h12;
      17'd39603: data = 8'h02;
      17'd39604: data = 8'hf4;
      17'd39605: data = 8'hfc;
      17'd39606: data = 8'hf2;
      17'd39607: data = 8'h15;
      17'd39608: data = 8'h0c;
      17'd39609: data = 8'hf4;
      17'd39610: data = 8'hf6;
      17'd39611: data = 8'hfc;
      17'd39612: data = 8'h0a;
      17'd39613: data = 8'h09;
      17'd39614: data = 8'h06;
      17'd39615: data = 8'hf2;
      17'd39616: data = 8'hef;
      17'd39617: data = 8'h06;
      17'd39618: data = 8'h16;
      17'd39619: data = 8'h09;
      17'd39620: data = 8'hda;
      17'd39621: data = 8'hf5;
      17'd39622: data = 8'h1b;
      17'd39623: data = 8'h09;
      17'd39624: data = 8'h09;
      17'd39625: data = 8'he2;
      17'd39626: data = 8'heb;
      17'd39627: data = 8'h24;
      17'd39628: data = 8'h0c;
      17'd39629: data = 8'hf9;
      17'd39630: data = 8'he2;
      17'd39631: data = 8'hf2;
      17'd39632: data = 8'h1e;
      17'd39633: data = 8'h13;
      17'd39634: data = 8'hf1;
      17'd39635: data = 8'he5;
      17'd39636: data = 8'h00;
      17'd39637: data = 8'h0c;
      17'd39638: data = 8'h06;
      17'd39639: data = 8'h05;
      17'd39640: data = 8'h0a;
      17'd39641: data = 8'hf1;
      17'd39642: data = 8'hf2;
      17'd39643: data = 8'h22;
      17'd39644: data = 8'hfc;
      17'd39645: data = 8'h02;
      17'd39646: data = 8'h0a;
      17'd39647: data = 8'he7;
      17'd39648: data = 8'h15;
      17'd39649: data = 8'h04;
      17'd39650: data = 8'hf6;
      17'd39651: data = 8'h11;
      17'd39652: data = 8'h04;
      17'd39653: data = 8'hf9;
      17'd39654: data = 8'hfd;
      17'd39655: data = 8'hfd;
      17'd39656: data = 8'h12;
      17'd39657: data = 8'h04;
      17'd39658: data = 8'he9;
      17'd39659: data = 8'h05;
      17'd39660: data = 8'h11;
      17'd39661: data = 8'h01;
      17'd39662: data = 8'hf4;
      17'd39663: data = 8'h06;
      17'd39664: data = 8'hfe;
      17'd39665: data = 8'hf6;
      17'd39666: data = 8'h12;
      17'd39667: data = 8'h00;
      17'd39668: data = 8'hf4;
      17'd39669: data = 8'h06;
      17'd39670: data = 8'h02;
      17'd39671: data = 8'h01;
      17'd39672: data = 8'h02;
      17'd39673: data = 8'h00;
      17'd39674: data = 8'h02;
      17'd39675: data = 8'hf6;
      17'd39676: data = 8'h0c;
      17'd39677: data = 8'h11;
      17'd39678: data = 8'hec;
      17'd39679: data = 8'hfa;
      17'd39680: data = 8'h13;
      17'd39681: data = 8'h0a;
      17'd39682: data = 8'he5;
      17'd39683: data = 8'hf9;
      17'd39684: data = 8'h1e;
      17'd39685: data = 8'hf6;
      17'd39686: data = 8'hfe;
      17'd39687: data = 8'h01;
      17'd39688: data = 8'hf2;
      17'd39689: data = 8'h0e;
      17'd39690: data = 8'h04;
      17'd39691: data = 8'hfa;
      17'd39692: data = 8'hf5;
      17'd39693: data = 8'h00;
      17'd39694: data = 8'hfd;
      17'd39695: data = 8'hf6;
      17'd39696: data = 8'h12;
      17'd39697: data = 8'h09;
      17'd39698: data = 8'hde;
      17'd39699: data = 8'hf4;
      17'd39700: data = 8'h1a;
      17'd39701: data = 8'h0a;
      17'd39702: data = 8'hfc;
      17'd39703: data = 8'he9;
      17'd39704: data = 8'hed;
      17'd39705: data = 8'h0c;
      17'd39706: data = 8'h2b;
      17'd39707: data = 8'h02;
      17'd39708: data = 8'hc6;
      17'd39709: data = 8'hf6;
      17'd39710: data = 8'h19;
      17'd39711: data = 8'h0a;
      17'd39712: data = 8'h1a;
      17'd39713: data = 8'hf2;
      17'd39714: data = 8'hc4;
      17'd39715: data = 8'h0d;
      17'd39716: data = 8'h31;
      17'd39717: data = 8'h04;
      17'd39718: data = 8'hf5;
      17'd39719: data = 8'hda;
      17'd39720: data = 8'hf4;
      17'd39721: data = 8'h2b;
      17'd39722: data = 8'h12;
      17'd39723: data = 8'hf6;
      17'd39724: data = 8'hdc;
      17'd39725: data = 8'hf9;
      17'd39726: data = 8'h26;
      17'd39727: data = 8'h06;
      17'd39728: data = 8'hed;
      17'd39729: data = 8'hfd;
      17'd39730: data = 8'hf5;
      17'd39731: data = 8'h09;
      17'd39732: data = 8'h1e;
      17'd39733: data = 8'heb;
      17'd39734: data = 8'hec;
      17'd39735: data = 8'h09;
      17'd39736: data = 8'h0e;
      17'd39737: data = 8'h02;
      17'd39738: data = 8'he9;
      17'd39739: data = 8'hf6;
      17'd39740: data = 8'h09;
      17'd39741: data = 8'h0d;
      17'd39742: data = 8'h06;
      17'd39743: data = 8'he9;
      17'd39744: data = 8'hf6;
      17'd39745: data = 8'h12;
      17'd39746: data = 8'hf6;
      17'd39747: data = 8'h0a;
      17'd39748: data = 8'h0d;
      17'd39749: data = 8'he2;
      17'd39750: data = 8'hf5;
      17'd39751: data = 8'h13;
      17'd39752: data = 8'h01;
      17'd39753: data = 8'h00;
      17'd39754: data = 8'hf4;
      17'd39755: data = 8'heb;
      17'd39756: data = 8'h13;
      17'd39757: data = 8'hfa;
      17'd39758: data = 8'hf5;
      17'd39759: data = 8'h0c;
      17'd39760: data = 8'hfe;
      17'd39761: data = 8'h02;
      17'd39762: data = 8'he7;
      17'd39763: data = 8'hfe;
      17'd39764: data = 8'h12;
      17'd39765: data = 8'hf9;
      17'd39766: data = 8'hf6;
      17'd39767: data = 8'h05;
      17'd39768: data = 8'hed;
      17'd39769: data = 8'hf6;
      17'd39770: data = 8'h23;
      17'd39771: data = 8'hef;
      17'd39772: data = 8'hf6;
      17'd39773: data = 8'hfc;
      17'd39774: data = 8'h05;
      17'd39775: data = 8'h0d;
      17'd39776: data = 8'hdc;
      17'd39777: data = 8'h09;
      17'd39778: data = 8'h13;
      17'd39779: data = 8'hf1;
      17'd39780: data = 8'h04;
      17'd39781: data = 8'h00;
      17'd39782: data = 8'he2;
      17'd39783: data = 8'h01;
      17'd39784: data = 8'h26;
      17'd39785: data = 8'hf9;
      17'd39786: data = 8'he5;
      17'd39787: data = 8'h02;
      17'd39788: data = 8'hf6;
      17'd39789: data = 8'h13;
      17'd39790: data = 8'h13;
      17'd39791: data = 8'hde;
      17'd39792: data = 8'hef;
      17'd39793: data = 8'hfc;
      17'd39794: data = 8'h0c;
      17'd39795: data = 8'h1a;
      17'd39796: data = 8'he4;
      17'd39797: data = 8'hdc;
      17'd39798: data = 8'h02;
      17'd39799: data = 8'h19;
      17'd39800: data = 8'h04;
      17'd39801: data = 8'hed;
      17'd39802: data = 8'heb;
      17'd39803: data = 8'h06;
      17'd39804: data = 8'h0e;
      17'd39805: data = 8'hfc;
      17'd39806: data = 8'h01;
      17'd39807: data = 8'hf2;
      17'd39808: data = 8'hfd;
      17'd39809: data = 8'h0c;
      17'd39810: data = 8'hfe;
      17'd39811: data = 8'hec;
      17'd39812: data = 8'hf5;
      17'd39813: data = 8'h0d;
      17'd39814: data = 8'h09;
      17'd39815: data = 8'hfd;
      17'd39816: data = 8'hed;
      17'd39817: data = 8'hf4;
      17'd39818: data = 8'h15;
      17'd39819: data = 8'hf6;
      17'd39820: data = 8'hfd;
      17'd39821: data = 8'h15;
      17'd39822: data = 8'hed;
      17'd39823: data = 8'h00;
      17'd39824: data = 8'h06;
      17'd39825: data = 8'hf2;
      17'd39826: data = 8'h09;
      17'd39827: data = 8'h15;
      17'd39828: data = 8'hf9;
      17'd39829: data = 8'hdc;
      17'd39830: data = 8'h01;
      17'd39831: data = 8'h19;
      17'd39832: data = 8'h0c;
      17'd39833: data = 8'hfe;
      17'd39834: data = 8'heb;
      17'd39835: data = 8'hec;
      17'd39836: data = 8'h06;
      17'd39837: data = 8'h11;
      17'd39838: data = 8'hfc;
      17'd39839: data = 8'h00;
      17'd39840: data = 8'he7;
      17'd39841: data = 8'hec;
      17'd39842: data = 8'h1b;
      17'd39843: data = 8'h01;
      17'd39844: data = 8'hfe;
      17'd39845: data = 8'hf6;
      17'd39846: data = 8'he5;
      17'd39847: data = 8'h04;
      17'd39848: data = 8'h0c;
      17'd39849: data = 8'h06;
      17'd39850: data = 8'hf4;
      17'd39851: data = 8'hf9;
      17'd39852: data = 8'hfc;
      17'd39853: data = 8'hfc;
      17'd39854: data = 8'h0d;
      17'd39855: data = 8'hfa;
      17'd39856: data = 8'hf5;
      17'd39857: data = 8'hfe;
      17'd39858: data = 8'hf1;
      17'd39859: data = 8'h04;
      17'd39860: data = 8'h0d;
      17'd39861: data = 8'hf6;
      17'd39862: data = 8'hfa;
      17'd39863: data = 8'h02;
      17'd39864: data = 8'hf6;
      17'd39865: data = 8'hfd;
      17'd39866: data = 8'h04;
      17'd39867: data = 8'hfd;
      17'd39868: data = 8'h0a;
      17'd39869: data = 8'hfc;
      17'd39870: data = 8'hf5;
      17'd39871: data = 8'h05;
      17'd39872: data = 8'hfc;
      17'd39873: data = 8'h04;
      17'd39874: data = 8'h02;
      17'd39875: data = 8'hfc;
      17'd39876: data = 8'h01;
      17'd39877: data = 8'h09;
      17'd39878: data = 8'h00;
      17'd39879: data = 8'hfe;
      17'd39880: data = 8'h02;
      17'd39881: data = 8'h01;
      17'd39882: data = 8'h0c;
      17'd39883: data = 8'h04;
      17'd39884: data = 8'hef;
      17'd39885: data = 8'h04;
      17'd39886: data = 8'h05;
      17'd39887: data = 8'h05;
      17'd39888: data = 8'h15;
      17'd39889: data = 8'he9;
      17'd39890: data = 8'hef;
      17'd39891: data = 8'h09;
      17'd39892: data = 8'h0c;
      17'd39893: data = 8'h05;
      17'd39894: data = 8'hed;
      17'd39895: data = 8'hfc;
      17'd39896: data = 8'h05;
      17'd39897: data = 8'hfc;
      17'd39898: data = 8'h05;
      17'd39899: data = 8'h00;
      17'd39900: data = 8'heb;
      17'd39901: data = 8'h06;
      17'd39902: data = 8'h0d;
      17'd39903: data = 8'hf9;
      17'd39904: data = 8'hfd;
      17'd39905: data = 8'h01;
      17'd39906: data = 8'h13;
      17'd39907: data = 8'hf9;
      17'd39908: data = 8'hec;
      17'd39909: data = 8'h0c;
      17'd39910: data = 8'h05;
      17'd39911: data = 8'h05;
      17'd39912: data = 8'hfc;
      17'd39913: data = 8'heb;
      17'd39914: data = 8'hfd;
      17'd39915: data = 8'h1c;
      17'd39916: data = 8'h06;
      17'd39917: data = 8'he4;
      17'd39918: data = 8'hfd;
      17'd39919: data = 8'h00;
      17'd39920: data = 8'hfe;
      17'd39921: data = 8'h0e;
      17'd39922: data = 8'h00;
      17'd39923: data = 8'hf4;
      17'd39924: data = 8'h02;
      17'd39925: data = 8'h00;
      17'd39926: data = 8'h04;
      17'd39927: data = 8'hfe;
      17'd39928: data = 8'hf5;
      17'd39929: data = 8'h13;
      17'd39930: data = 8'hfd;
      17'd39931: data = 8'hf9;
      17'd39932: data = 8'h0d;
      17'd39933: data = 8'hec;
      17'd39934: data = 8'h05;
      17'd39935: data = 8'h1f;
      17'd39936: data = 8'he9;
      17'd39937: data = 8'heb;
      17'd39938: data = 8'h0a;
      17'd39939: data = 8'h09;
      17'd39940: data = 8'h06;
      17'd39941: data = 8'h01;
      17'd39942: data = 8'heb;
      17'd39943: data = 8'hf5;
      17'd39944: data = 8'h19;
      17'd39945: data = 8'h05;
      17'd39946: data = 8'hed;
      17'd39947: data = 8'hf4;
      17'd39948: data = 8'hfe;
      17'd39949: data = 8'h13;
      17'd39950: data = 8'h05;
      17'd39951: data = 8'hf6;
      17'd39952: data = 8'hf1;
      17'd39953: data = 8'h00;
      17'd39954: data = 8'h0d;
      17'd39955: data = 8'h00;
      17'd39956: data = 8'hf9;
      17'd39957: data = 8'hf4;
      17'd39958: data = 8'h04;
      17'd39959: data = 8'h0d;
      17'd39960: data = 8'h02;
      17'd39961: data = 8'hed;
      17'd39962: data = 8'hfa;
      17'd39963: data = 8'h0d;
      17'd39964: data = 8'h04;
      17'd39965: data = 8'h02;
      17'd39966: data = 8'hf9;
      17'd39967: data = 8'hfa;
      17'd39968: data = 8'h0a;
      17'd39969: data = 8'h0c;
      17'd39970: data = 8'hfd;
      17'd39971: data = 8'hf1;
      17'd39972: data = 8'h00;
      17'd39973: data = 8'h06;
      17'd39974: data = 8'h05;
      17'd39975: data = 8'hfd;
      17'd39976: data = 8'h00;
      17'd39977: data = 8'h02;
      17'd39978: data = 8'h01;
      17'd39979: data = 8'h00;
      17'd39980: data = 8'hfe;
      17'd39981: data = 8'h06;
      17'd39982: data = 8'hf6;
      17'd39983: data = 8'h00;
      17'd39984: data = 8'h04;
      17'd39985: data = 8'hfc;
      17'd39986: data = 8'h01;
      17'd39987: data = 8'hfa;
      17'd39988: data = 8'hfd;
      17'd39989: data = 8'h00;
      17'd39990: data = 8'hf9;
      17'd39991: data = 8'hfa;
      17'd39992: data = 8'h01;
      17'd39993: data = 8'h00;
      17'd39994: data = 8'hfd;
      17'd39995: data = 8'hfa;
      17'd39996: data = 8'hfe;
      17'd39997: data = 8'h06;
      17'd39998: data = 8'h00;
      17'd39999: data = 8'hed;
      17'd40000: data = 8'hfa;
      17'd40001: data = 8'h06;
      17'd40002: data = 8'h01;
      17'd40003: data = 8'h01;
      17'd40004: data = 8'hfc;
      17'd40005: data = 8'hfc;
      17'd40006: data = 8'h00;
      17'd40007: data = 8'h0a;
      17'd40008: data = 8'h02;
      17'd40009: data = 8'hf5;
      17'd40010: data = 8'hfe;
      17'd40011: data = 8'h04;
      17'd40012: data = 8'h09;
      17'd40013: data = 8'hfc;
      17'd40014: data = 8'hfa;
      17'd40015: data = 8'h04;
      17'd40016: data = 8'h04;
      17'd40017: data = 8'h04;
      17'd40018: data = 8'hf4;
      17'd40019: data = 8'h01;
      17'd40020: data = 8'h0d;
      17'd40021: data = 8'hf9;
      17'd40022: data = 8'h01;
      17'd40023: data = 8'h04;
      17'd40024: data = 8'hfe;
      17'd40025: data = 8'h02;
      17'd40026: data = 8'h05;
      17'd40027: data = 8'hfd;
      17'd40028: data = 8'hf9;
      17'd40029: data = 8'h01;
      17'd40030: data = 8'h09;
      17'd40031: data = 8'h04;
      17'd40032: data = 8'hf9;
      17'd40033: data = 8'hfa;
      17'd40034: data = 8'h00;
      17'd40035: data = 8'h01;
      17'd40036: data = 8'h0a;
      17'd40037: data = 8'hfc;
      17'd40038: data = 8'hf2;
      17'd40039: data = 8'h01;
      17'd40040: data = 8'h05;
      17'd40041: data = 8'h04;
      17'd40042: data = 8'hfc;
      17'd40043: data = 8'hf9;
      17'd40044: data = 8'hfc;
      17'd40045: data = 8'h05;
      17'd40046: data = 8'h05;
      17'd40047: data = 8'hf6;
      17'd40048: data = 8'hfa;
      17'd40049: data = 8'hfa;
      17'd40050: data = 8'h01;
      17'd40051: data = 8'h02;
      17'd40052: data = 8'hfe;
      17'd40053: data = 8'h01;
      17'd40054: data = 8'hf1;
      17'd40055: data = 8'h00;
      17'd40056: data = 8'h00;
      17'd40057: data = 8'hf4;
      17'd40058: data = 8'h09;
      17'd40059: data = 8'h04;
      17'd40060: data = 8'hf4;
      17'd40061: data = 8'hfd;
      17'd40062: data = 8'h00;
      17'd40063: data = 8'h01;
      17'd40064: data = 8'h06;
      17'd40065: data = 8'hf6;
      17'd40066: data = 8'h01;
      17'd40067: data = 8'h00;
      17'd40068: data = 8'hf9;
      17'd40069: data = 8'h09;
      17'd40070: data = 8'hfa;
      17'd40071: data = 8'hfd;
      17'd40072: data = 8'h09;
      17'd40073: data = 8'hfd;
      17'd40074: data = 8'hf9;
      17'd40075: data = 8'h01;
      17'd40076: data = 8'h01;
      17'd40077: data = 8'h00;
      17'd40078: data = 8'hfe;
      17'd40079: data = 8'hf6;
      17'd40080: data = 8'h02;
      17'd40081: data = 8'h0c;
      17'd40082: data = 8'hf9;
      17'd40083: data = 8'hf6;
      17'd40084: data = 8'h01;
      17'd40085: data = 8'hfc;
      17'd40086: data = 8'h02;
      17'd40087: data = 8'h05;
      17'd40088: data = 8'hfa;
      17'd40089: data = 8'hfa;
      17'd40090: data = 8'hfa;
      17'd40091: data = 8'h06;
      17'd40092: data = 8'h09;
      17'd40093: data = 8'hfa;
      17'd40094: data = 8'hfc;
      17'd40095: data = 8'hf5;
      17'd40096: data = 8'hfe;
      17'd40097: data = 8'h0d;
      17'd40098: data = 8'hfd;
      17'd40099: data = 8'hf6;
      17'd40100: data = 8'hfd;
      17'd40101: data = 8'h01;
      17'd40102: data = 8'h00;
      17'd40103: data = 8'hfd;
      17'd40104: data = 8'hfd;
      17'd40105: data = 8'hfa;
      17'd40106: data = 8'h01;
      17'd40107: data = 8'h01;
      17'd40108: data = 8'h00;
      17'd40109: data = 8'h04;
      17'd40110: data = 8'h00;
      17'd40111: data = 8'hfd;
      17'd40112: data = 8'h02;
      17'd40113: data = 8'h02;
      17'd40114: data = 8'hfd;
      17'd40115: data = 8'h00;
      17'd40116: data = 8'h01;
      17'd40117: data = 8'h00;
      17'd40118: data = 8'hfe;
      17'd40119: data = 8'h02;
      17'd40120: data = 8'h02;
      17'd40121: data = 8'hfd;
      17'd40122: data = 8'hfe;
      17'd40123: data = 8'h01;
      17'd40124: data = 8'hfc;
      17'd40125: data = 8'h09;
      17'd40126: data = 8'h05;
      17'd40127: data = 8'hf4;
      17'd40128: data = 8'hfe;
      17'd40129: data = 8'h05;
      17'd40130: data = 8'h01;
      17'd40131: data = 8'h02;
      17'd40132: data = 8'hfe;
      17'd40133: data = 8'hf6;
      17'd40134: data = 8'h02;
      17'd40135: data = 8'h06;
      17'd40136: data = 8'hfe;
      17'd40137: data = 8'h04;
      17'd40138: data = 8'h02;
      17'd40139: data = 8'hfc;
      17'd40140: data = 8'h02;
      17'd40141: data = 8'h01;
      17'd40142: data = 8'hfe;
      17'd40143: data = 8'h04;
      17'd40144: data = 8'h00;
      17'd40145: data = 8'hfd;
      17'd40146: data = 8'h02;
      17'd40147: data = 8'h01;
      17'd40148: data = 8'h01;
      17'd40149: data = 8'h00;
      17'd40150: data = 8'hfc;
      17'd40151: data = 8'hfe;
      17'd40152: data = 8'h02;
      17'd40153: data = 8'h05;
      17'd40154: data = 8'h04;
      17'd40155: data = 8'hfc;
      17'd40156: data = 8'hfc;
      17'd40157: data = 8'h01;
      17'd40158: data = 8'h02;
      17'd40159: data = 8'h01;
      17'd40160: data = 8'h00;
      17'd40161: data = 8'hfd;
      17'd40162: data = 8'hfe;
      17'd40163: data = 8'h02;
      17'd40164: data = 8'h04;
      17'd40165: data = 8'h04;
      17'd40166: data = 8'h00;
      17'd40167: data = 8'hf9;
      17'd40168: data = 8'h00;
      17'd40169: data = 8'h04;
      17'd40170: data = 8'h04;
      17'd40171: data = 8'h02;
      17'd40172: data = 8'hfc;
      17'd40173: data = 8'hfe;
      17'd40174: data = 8'h00;
      17'd40175: data = 8'h01;
      17'd40176: data = 8'h00;
      17'd40177: data = 8'hfa;
      17'd40178: data = 8'hf9;
      17'd40179: data = 8'hfe;
      17'd40180: data = 8'h04;
      17'd40181: data = 8'hfe;
      17'd40182: data = 8'hfa;
      17'd40183: data = 8'hfc;
      17'd40184: data = 8'h00;
      17'd40185: data = 8'h00;
      17'd40186: data = 8'h00;
      17'd40187: data = 8'hfa;
      17'd40188: data = 8'hf9;
      17'd40189: data = 8'h01;
      17'd40190: data = 8'h02;
      17'd40191: data = 8'h00;
      17'd40192: data = 8'hfc;
      17'd40193: data = 8'hfc;
      17'd40194: data = 8'hfe;
      17'd40195: data = 8'hfd;
      17'd40196: data = 8'hfd;
      17'd40197: data = 8'hfe;
      17'd40198: data = 8'hfe;
      17'd40199: data = 8'h00;
      17'd40200: data = 8'h02;
      17'd40201: data = 8'hfd;
      17'd40202: data = 8'hf6;
      17'd40203: data = 8'h01;
      17'd40204: data = 8'h04;
      17'd40205: data = 8'h00;
      17'd40206: data = 8'hfd;
      17'd40207: data = 8'hfa;
      17'd40208: data = 8'h04;
      17'd40209: data = 8'h04;
      17'd40210: data = 8'hfe;
      17'd40211: data = 8'h01;
      17'd40212: data = 8'hfd;
      17'd40213: data = 8'h00;
      17'd40214: data = 8'h02;
      17'd40215: data = 8'hfd;
      17'd40216: data = 8'h02;
      17'd40217: data = 8'h00;
      17'd40218: data = 8'hfa;
      17'd40219: data = 8'h01;
      17'd40220: data = 8'h01;
      17'd40221: data = 8'hfe;
      17'd40222: data = 8'hfd;
      17'd40223: data = 8'hfd;
      17'd40224: data = 8'hfc;
      17'd40225: data = 8'h02;
      17'd40226: data = 8'h00;
      17'd40227: data = 8'hfd;
      17'd40228: data = 8'h01;
      17'd40229: data = 8'h00;
      17'd40230: data = 8'hfd;
      17'd40231: data = 8'hfd;
      17'd40232: data = 8'hfe;
      17'd40233: data = 8'h02;
      17'd40234: data = 8'h02;
      17'd40235: data = 8'hfd;
      17'd40236: data = 8'hfd;
      17'd40237: data = 8'hfe;
      17'd40238: data = 8'h00;
      17'd40239: data = 8'hfe;
      17'd40240: data = 8'hfd;
      17'd40241: data = 8'hfe;
      17'd40242: data = 8'hfd;
      17'd40243: data = 8'h01;
      17'd40244: data = 8'h00;
      17'd40245: data = 8'hfc;
      17'd40246: data = 8'h01;
      17'd40247: data = 8'h01;
      17'd40248: data = 8'h00;
      17'd40249: data = 8'h02;
      17'd40250: data = 8'hfd;
      17'd40251: data = 8'hfe;
      17'd40252: data = 8'h02;
      17'd40253: data = 8'hfe;
      17'd40254: data = 8'hfe;
      17'd40255: data = 8'hfe;
      17'd40256: data = 8'hfe;
      17'd40257: data = 8'h00;
      17'd40258: data = 8'h04;
      17'd40259: data = 8'h00;
      17'd40260: data = 8'hfc;
      17'd40261: data = 8'h02;
      17'd40262: data = 8'h04;
      17'd40263: data = 8'h04;
      17'd40264: data = 8'h09;
      17'd40265: data = 8'hfd;
      17'd40266: data = 8'hfe;
      17'd40267: data = 8'h04;
      17'd40268: data = 8'h04;
      17'd40269: data = 8'h05;
      17'd40270: data = 8'hfd;
      17'd40271: data = 8'hfd;
      17'd40272: data = 8'h00;
      17'd40273: data = 8'h04;
      17'd40274: data = 8'h01;
      17'd40275: data = 8'hfd;
      17'd40276: data = 8'hfe;
      17'd40277: data = 8'h01;
      17'd40278: data = 8'h01;
      17'd40279: data = 8'hfa;
      17'd40280: data = 8'h00;
      17'd40281: data = 8'h05;
      17'd40282: data = 8'hfe;
      17'd40283: data = 8'hfe;
      17'd40284: data = 8'hf9;
      17'd40285: data = 8'hfa;
      17'd40286: data = 8'h04;
      17'd40287: data = 8'h01;
      17'd40288: data = 8'hfd;
      17'd40289: data = 8'hf9;
      17'd40290: data = 8'hf9;
      17'd40291: data = 8'h01;
      17'd40292: data = 8'h04;
      17'd40293: data = 8'hfe;
      17'd40294: data = 8'hfa;
      17'd40295: data = 8'hf6;
      17'd40296: data = 8'h00;
      17'd40297: data = 8'hfe;
      17'd40298: data = 8'hfa;
      17'd40299: data = 8'h01;
      17'd40300: data = 8'hfc;
      17'd40301: data = 8'h00;
      17'd40302: data = 8'h01;
      17'd40303: data = 8'hfa;
      17'd40304: data = 8'hfe;
      17'd40305: data = 8'h00;
      17'd40306: data = 8'h04;
      17'd40307: data = 8'h02;
      17'd40308: data = 8'hfc;
      17'd40309: data = 8'hfc;
      17'd40310: data = 8'h00;
      17'd40311: data = 8'h02;
      17'd40312: data = 8'h04;
      17'd40313: data = 8'hfd;
      17'd40314: data = 8'hfc;
      17'd40315: data = 8'h01;
      17'd40316: data = 8'h00;
      17'd40317: data = 8'h01;
      17'd40318: data = 8'h00;
      17'd40319: data = 8'h00;
      17'd40320: data = 8'h00;
      17'd40321: data = 8'h01;
      17'd40322: data = 8'h01;
      17'd40323: data = 8'hfe;
      17'd40324: data = 8'h01;
      17'd40325: data = 8'h00;
      17'd40326: data = 8'h01;
      17'd40327: data = 8'h01;
      17'd40328: data = 8'hfe;
      17'd40329: data = 8'h00;
      17'd40330: data = 8'h00;
      17'd40331: data = 8'hfe;
      17'd40332: data = 8'hfe;
      17'd40333: data = 8'hfc;
      17'd40334: data = 8'hfe;
      17'd40335: data = 8'h02;
      17'd40336: data = 8'h00;
      17'd40337: data = 8'hfe;
      17'd40338: data = 8'hfd;
      17'd40339: data = 8'h01;
      17'd40340: data = 8'h01;
      17'd40341: data = 8'h01;
      17'd40342: data = 8'hfe;
      17'd40343: data = 8'hfc;
      17'd40344: data = 8'hfc;
      17'd40345: data = 8'hfd;
      17'd40346: data = 8'h00;
      17'd40347: data = 8'hfd;
      17'd40348: data = 8'hfa;
      17'd40349: data = 8'hfc;
      17'd40350: data = 8'hfd;
      17'd40351: data = 8'hfc;
      17'd40352: data = 8'hfe;
      17'd40353: data = 8'h01;
      17'd40354: data = 8'hfe;
      17'd40355: data = 8'h02;
      17'd40356: data = 8'h05;
      17'd40357: data = 8'h01;
      17'd40358: data = 8'hfe;
      17'd40359: data = 8'h02;
      17'd40360: data = 8'h04;
      17'd40361: data = 8'h04;
      17'd40362: data = 8'h01;
      17'd40363: data = 8'h00;
      17'd40364: data = 8'h04;
      17'd40365: data = 8'h04;
      17'd40366: data = 8'h05;
      17'd40367: data = 8'h05;
      17'd40368: data = 8'h01;
      17'd40369: data = 8'h02;
      17'd40370: data = 8'h04;
      17'd40371: data = 8'h02;
      17'd40372: data = 8'h04;
      17'd40373: data = 8'h00;
      17'd40374: data = 8'h04;
      17'd40375: data = 8'h05;
      17'd40376: data = 8'hfe;
      17'd40377: data = 8'h01;
      17'd40378: data = 8'h01;
      17'd40379: data = 8'hfe;
      17'd40380: data = 8'hfe;
      17'd40381: data = 8'h01;
      17'd40382: data = 8'h02;
      17'd40383: data = 8'h00;
      17'd40384: data = 8'h01;
      17'd40385: data = 8'h02;
      17'd40386: data = 8'hfe;
      17'd40387: data = 8'hfe;
      17'd40388: data = 8'h00;
      17'd40389: data = 8'hfa;
      17'd40390: data = 8'hfc;
      17'd40391: data = 8'hfe;
      17'd40392: data = 8'hf9;
      17'd40393: data = 8'hfa;
      17'd40394: data = 8'hfc;
      17'd40395: data = 8'hfc;
      17'd40396: data = 8'hf9;
      17'd40397: data = 8'hfa;
      17'd40398: data = 8'hf9;
      17'd40399: data = 8'hf6;
      17'd40400: data = 8'hf9;
      17'd40401: data = 8'hfa;
      17'd40402: data = 8'hfc;
      17'd40403: data = 8'hf9;
      17'd40404: data = 8'hfc;
      17'd40405: data = 8'hfa;
      17'd40406: data = 8'hf4;
      17'd40407: data = 8'hfc;
      17'd40408: data = 8'hfe;
      17'd40409: data = 8'hfc;
      17'd40410: data = 8'h02;
      17'd40411: data = 8'h01;
      17'd40412: data = 8'hfa;
      17'd40413: data = 8'h05;
      17'd40414: data = 8'h04;
      17'd40415: data = 8'h01;
      17'd40416: data = 8'h09;
      17'd40417: data = 8'h06;
      17'd40418: data = 8'h09;
      17'd40419: data = 8'h0a;
      17'd40420: data = 8'h0c;
      17'd40421: data = 8'h0d;
      17'd40422: data = 8'h0e;
      17'd40423: data = 8'h0c;
      17'd40424: data = 8'h0c;
      17'd40425: data = 8'h0e;
      17'd40426: data = 8'h0c;
      17'd40427: data = 8'h11;
      17'd40428: data = 8'h11;
      17'd40429: data = 8'h0a;
      17'd40430: data = 8'h09;
      17'd40431: data = 8'h0d;
      17'd40432: data = 8'h0a;
      17'd40433: data = 8'h09;
      17'd40434: data = 8'h0d;
      17'd40435: data = 8'h05;
      17'd40436: data = 8'h04;
      17'd40437: data = 8'h09;
      17'd40438: data = 8'h06;
      17'd40439: data = 8'h02;
      17'd40440: data = 8'h00;
      17'd40441: data = 8'hfe;
      17'd40442: data = 8'hfa;
      17'd40443: data = 8'hfa;
      17'd40444: data = 8'hfe;
      17'd40445: data = 8'hfa;
      17'd40446: data = 8'hf5;
      17'd40447: data = 8'hf5;
      17'd40448: data = 8'hf2;
      17'd40449: data = 8'hf9;
      17'd40450: data = 8'hf6;
      17'd40451: data = 8'hef;
      17'd40452: data = 8'hed;
      17'd40453: data = 8'hf2;
      17'd40454: data = 8'hf4;
      17'd40455: data = 8'hf2;
      17'd40456: data = 8'hef;
      17'd40457: data = 8'hed;
      17'd40458: data = 8'hef;
      17'd40459: data = 8'hf2;
      17'd40460: data = 8'hef;
      17'd40461: data = 8'hef;
      17'd40462: data = 8'hf4;
      17'd40463: data = 8'hf4;
      17'd40464: data = 8'hf6;
      17'd40465: data = 8'hf6;
      17'd40466: data = 8'hf2;
      17'd40467: data = 8'hf6;
      17'd40468: data = 8'hfc;
      17'd40469: data = 8'hf9;
      17'd40470: data = 8'hfa;
      17'd40471: data = 8'hfc;
      17'd40472: data = 8'hfc;
      17'd40473: data = 8'hfd;
      17'd40474: data = 8'hfe;
      17'd40475: data = 8'hfe;
      17'd40476: data = 8'h00;
      17'd40477: data = 8'hfe;
      17'd40478: data = 8'h00;
      17'd40479: data = 8'hfd;
      17'd40480: data = 8'h01;
      17'd40481: data = 8'h05;
      17'd40482: data = 8'h02;
      17'd40483: data = 8'h01;
      17'd40484: data = 8'h02;
      17'd40485: data = 8'h02;
      17'd40486: data = 8'h04;
      17'd40487: data = 8'h05;
      17'd40488: data = 8'hfe;
      17'd40489: data = 8'h01;
      17'd40490: data = 8'h01;
      17'd40491: data = 8'h01;
      17'd40492: data = 8'h06;
      17'd40493: data = 8'h00;
      17'd40494: data = 8'hfd;
      17'd40495: data = 8'h00;
      17'd40496: data = 8'h01;
      17'd40497: data = 8'hfe;
      17'd40498: data = 8'h00;
      17'd40499: data = 8'hfd;
      17'd40500: data = 8'hfc;
      17'd40501: data = 8'h04;
      17'd40502: data = 8'h02;
      17'd40503: data = 8'hfc;
      17'd40504: data = 8'hfd;
      17'd40505: data = 8'hfe;
      17'd40506: data = 8'hfc;
      17'd40507: data = 8'hfd;
      17'd40508: data = 8'hfc;
      17'd40509: data = 8'hf6;
      17'd40510: data = 8'hfa;
      17'd40511: data = 8'hfe;
      17'd40512: data = 8'h01;
      17'd40513: data = 8'hfd;
      17'd40514: data = 8'hfa;
      17'd40515: data = 8'hf9;
      17'd40516: data = 8'hfd;
      17'd40517: data = 8'h04;
      17'd40518: data = 8'h01;
      17'd40519: data = 8'h00;
      17'd40520: data = 8'hfd;
      17'd40521: data = 8'hfe;
      17'd40522: data = 8'h09;
      17'd40523: data = 8'h04;
      17'd40524: data = 8'h00;
      17'd40525: data = 8'h00;
      17'd40526: data = 8'hfe;
      17'd40527: data = 8'h04;
      17'd40528: data = 8'h0a;
      17'd40529: data = 8'h0a;
      17'd40530: data = 8'h02;
      17'd40531: data = 8'h01;
      17'd40532: data = 8'h0a;
      17'd40533: data = 8'h06;
      17'd40534: data = 8'h02;
      17'd40535: data = 8'h09;
      17'd40536: data = 8'hfe;
      17'd40537: data = 8'h00;
      17'd40538: data = 8'h09;
      17'd40539: data = 8'hfe;
      17'd40540: data = 8'h01;
      17'd40541: data = 8'h05;
      17'd40542: data = 8'h01;
      17'd40543: data = 8'h01;
      17'd40544: data = 8'hfe;
      17'd40545: data = 8'h01;
      17'd40546: data = 8'h04;
      17'd40547: data = 8'hfd;
      17'd40548: data = 8'h04;
      17'd40549: data = 8'h05;
      17'd40550: data = 8'hfa;
      17'd40551: data = 8'hfa;
      17'd40552: data = 8'hf6;
      17'd40553: data = 8'hf1;
      17'd40554: data = 8'hf6;
      17'd40555: data = 8'hfc;
      17'd40556: data = 8'hf9;
      17'd40557: data = 8'hf5;
      17'd40558: data = 8'hf6;
      17'd40559: data = 8'hfe;
      17'd40560: data = 8'h01;
      17'd40561: data = 8'hfd;
      17'd40562: data = 8'h01;
      17'd40563: data = 8'h04;
      17'd40564: data = 8'h04;
      17'd40565: data = 8'h09;
      17'd40566: data = 8'h0a;
      17'd40567: data = 8'h05;
      17'd40568: data = 8'h05;
      17'd40569: data = 8'h0d;
      17'd40570: data = 8'h0a;
      17'd40571: data = 8'h06;
      17'd40572: data = 8'h04;
      17'd40573: data = 8'h0a;
      17'd40574: data = 8'h0e;
      17'd40575: data = 8'h0a;
      17'd40576: data = 8'h13;
      17'd40577: data = 8'h0e;
      17'd40578: data = 8'h0a;
      17'd40579: data = 8'h11;
      17'd40580: data = 8'h0c;
      17'd40581: data = 8'h06;
      17'd40582: data = 8'h09;
      17'd40583: data = 8'h09;
      17'd40584: data = 8'h04;
      17'd40585: data = 8'h01;
      17'd40586: data = 8'h01;
      17'd40587: data = 8'hfc;
      17'd40588: data = 8'hf5;
      17'd40589: data = 8'hf9;
      17'd40590: data = 8'hfc;
      17'd40591: data = 8'hf9;
      17'd40592: data = 8'hf6;
      17'd40593: data = 8'hf4;
      17'd40594: data = 8'hf5;
      17'd40595: data = 8'hf9;
      17'd40596: data = 8'hf9;
      17'd40597: data = 8'hf5;
      17'd40598: data = 8'hed;
      17'd40599: data = 8'hed;
      17'd40600: data = 8'hf2;
      17'd40601: data = 8'hf1;
      17'd40602: data = 8'hec;
      17'd40603: data = 8'he7;
      17'd40604: data = 8'he9;
      17'd40605: data = 8'hec;
      17'd40606: data = 8'he9;
      17'd40607: data = 8'he9;
      17'd40608: data = 8'he9;
      17'd40609: data = 8'heb;
      17'd40610: data = 8'hf1;
      17'd40611: data = 8'hf2;
      17'd40612: data = 8'hf6;
      17'd40613: data = 8'hf9;
      17'd40614: data = 8'hfa;
      17'd40615: data = 8'hfd;
      17'd40616: data = 8'h01;
      17'd40617: data = 8'h02;
      17'd40618: data = 8'h01;
      17'd40619: data = 8'h06;
      17'd40620: data = 8'h09;
      17'd40621: data = 8'h0e;
      17'd40622: data = 8'h15;
      17'd40623: data = 8'h0d;
      17'd40624: data = 8'h12;
      17'd40625: data = 8'h1c;
      17'd40626: data = 8'h1b;
      17'd40627: data = 8'h1a;
      17'd40628: data = 8'h1a;
      17'd40629: data = 8'h1c;
      17'd40630: data = 8'h1f;
      17'd40631: data = 8'h22;
      17'd40632: data = 8'h22;
      17'd40633: data = 8'h1a;
      17'd40634: data = 8'h1a;
      17'd40635: data = 8'h1b;
      17'd40636: data = 8'h19;
      17'd40637: data = 8'h19;
      17'd40638: data = 8'h15;
      17'd40639: data = 8'h0d;
      17'd40640: data = 8'h0d;
      17'd40641: data = 8'h0c;
      17'd40642: data = 8'h0a;
      17'd40643: data = 8'h06;
      17'd40644: data = 8'hfe;
      17'd40645: data = 8'hfd;
      17'd40646: data = 8'hfd;
      17'd40647: data = 8'hfa;
      17'd40648: data = 8'hfa;
      17'd40649: data = 8'hf4;
      17'd40650: data = 8'hf1;
      17'd40651: data = 8'hef;
      17'd40652: data = 8'hed;
      17'd40653: data = 8'hed;
      17'd40654: data = 8'he9;
      17'd40655: data = 8'he9;
      17'd40656: data = 8'he5;
      17'd40657: data = 8'heb;
      17'd40658: data = 8'heb;
      17'd40659: data = 8'he9;
      17'd40660: data = 8'he9;
      17'd40661: data = 8'he7;
      17'd40662: data = 8'heb;
      17'd40663: data = 8'hed;
      17'd40664: data = 8'hed;
      17'd40665: data = 8'hef;
      17'd40666: data = 8'hf2;
      17'd40667: data = 8'hf5;
      17'd40668: data = 8'hf5;
      17'd40669: data = 8'hfa;
      17'd40670: data = 8'hfa;
      17'd40671: data = 8'hf5;
      17'd40672: data = 8'hfa;
      17'd40673: data = 8'hfe;
      17'd40674: data = 8'h01;
      17'd40675: data = 8'h05;
      17'd40676: data = 8'h05;
      17'd40677: data = 8'hfe;
      17'd40678: data = 8'h00;
      17'd40679: data = 8'h0a;
      17'd40680: data = 8'h06;
      17'd40681: data = 8'h05;
      17'd40682: data = 8'h02;
      17'd40683: data = 8'h01;
      17'd40684: data = 8'hfe;
      17'd40685: data = 8'h04;
      17'd40686: data = 8'h05;
      17'd40687: data = 8'hfc;
      17'd40688: data = 8'hfe;
      17'd40689: data = 8'hfe;
      17'd40690: data = 8'hfc;
      17'd40691: data = 8'hfa;
      17'd40692: data = 8'hfa;
      17'd40693: data = 8'hfc;
      17'd40694: data = 8'hf6;
      17'd40695: data = 8'hf6;
      17'd40696: data = 8'hf4;
      17'd40697: data = 8'hef;
      17'd40698: data = 8'hef;
      17'd40699: data = 8'hf1;
      17'd40700: data = 8'hef;
      17'd40701: data = 8'he9;
      17'd40702: data = 8'heb;
      17'd40703: data = 8'hf1;
      17'd40704: data = 8'heb;
      17'd40705: data = 8'hef;
      17'd40706: data = 8'hef;
      17'd40707: data = 8'he9;
      17'd40708: data = 8'heb;
      17'd40709: data = 8'hf1;
      17'd40710: data = 8'hed;
      17'd40711: data = 8'heb;
      17'd40712: data = 8'hf4;
      17'd40713: data = 8'hf1;
      17'd40714: data = 8'hf2;
      17'd40715: data = 8'hf4;
      17'd40716: data = 8'hf4;
      17'd40717: data = 8'hf5;
      17'd40718: data = 8'hf9;
      17'd40719: data = 8'hfe;
      17'd40720: data = 8'hfc;
      17'd40721: data = 8'h01;
      17'd40722: data = 8'h01;
      17'd40723: data = 8'h02;
      17'd40724: data = 8'h02;
      17'd40725: data = 8'h02;
      17'd40726: data = 8'h05;
      17'd40727: data = 8'h02;
      17'd40728: data = 8'h06;
      17'd40729: data = 8'h0a;
      17'd40730: data = 8'h09;
      17'd40731: data = 8'h0a;
      17'd40732: data = 8'h0a;
      17'd40733: data = 8'h0a;
      17'd40734: data = 8'h0e;
      17'd40735: data = 8'h0c;
      17'd40736: data = 8'h06;
      17'd40737: data = 8'h06;
      17'd40738: data = 8'h0d;
      17'd40739: data = 8'h0e;
      17'd40740: data = 8'h09;
      17'd40741: data = 8'h05;
      17'd40742: data = 8'h04;
      17'd40743: data = 8'h02;
      17'd40744: data = 8'h02;
      17'd40745: data = 8'h06;
      17'd40746: data = 8'h05;
      17'd40747: data = 8'h01;
      17'd40748: data = 8'h02;
      17'd40749: data = 8'h05;
      17'd40750: data = 8'h05;
      17'd40751: data = 8'h02;
      17'd40752: data = 8'h04;
      17'd40753: data = 8'h02;
      17'd40754: data = 8'h01;
      17'd40755: data = 8'h04;
      17'd40756: data = 8'h01;
      17'd40757: data = 8'hfe;
      17'd40758: data = 8'hfe;
      17'd40759: data = 8'h02;
      17'd40760: data = 8'h04;
      17'd40761: data = 8'hfd;
      17'd40762: data = 8'hfe;
      17'd40763: data = 8'h04;
      17'd40764: data = 8'h02;
      17'd40765: data = 8'h05;
      17'd40766: data = 8'h04;
      17'd40767: data = 8'h04;
      17'd40768: data = 8'h05;
      17'd40769: data = 8'h04;
      17'd40770: data = 8'h0a;
      17'd40771: data = 8'h06;
      17'd40772: data = 8'h05;
      17'd40773: data = 8'h05;
      17'd40774: data = 8'h05;
      17'd40775: data = 8'h0c;
      17'd40776: data = 8'h0e;
      17'd40777: data = 8'h13;
      17'd40778: data = 8'h0c;
      17'd40779: data = 8'h06;
      17'd40780: data = 8'h15;
      17'd40781: data = 8'h11;
      17'd40782: data = 8'h0d;
      17'd40783: data = 8'h12;
      17'd40784: data = 8'h0a;
      17'd40785: data = 8'h0d;
      17'd40786: data = 8'h0d;
      17'd40787: data = 8'h09;
      17'd40788: data = 8'h0a;
      17'd40789: data = 8'h05;
      17'd40790: data = 8'h09;
      17'd40791: data = 8'h0e;
      17'd40792: data = 8'h0c;
      17'd40793: data = 8'h0a;
      17'd40794: data = 8'h0e;
      17'd40795: data = 8'h0a;
      17'd40796: data = 8'h05;
      17'd40797: data = 8'h0a;
      17'd40798: data = 8'h02;
      17'd40799: data = 8'hf9;
      17'd40800: data = 8'hfd;
      17'd40801: data = 8'hfe;
      17'd40802: data = 8'hfe;
      17'd40803: data = 8'hfe;
      17'd40804: data = 8'hfa;
      17'd40805: data = 8'hfa;
      17'd40806: data = 8'hf9;
      17'd40807: data = 8'hfe;
      17'd40808: data = 8'h09;
      17'd40809: data = 8'hfd;
      17'd40810: data = 8'h00;
      17'd40811: data = 8'h12;
      17'd40812: data = 8'h0d;
      17'd40813: data = 8'h0e;
      17'd40814: data = 8'h12;
      17'd40815: data = 8'h12;
      17'd40816: data = 8'h11;
      17'd40817: data = 8'h11;
      17'd40818: data = 8'h13;
      17'd40819: data = 8'h0e;
      17'd40820: data = 8'h0d;
      17'd40821: data = 8'h12;
      17'd40822: data = 8'h13;
      17'd40823: data = 8'h0e;
      17'd40824: data = 8'h0d;
      17'd40825: data = 8'h0e;
      17'd40826: data = 8'h09;
      17'd40827: data = 8'h09;
      17'd40828: data = 8'h0e;
      17'd40829: data = 8'h06;
      17'd40830: data = 8'h02;
      17'd40831: data = 8'h09;
      17'd40832: data = 8'h01;
      17'd40833: data = 8'hfa;
      17'd40834: data = 8'hf6;
      17'd40835: data = 8'hf5;
      17'd40836: data = 8'hf2;
      17'd40837: data = 8'hed;
      17'd40838: data = 8'he9;
      17'd40839: data = 8'he5;
      17'd40840: data = 8'he5;
      17'd40841: data = 8'he4;
      17'd40842: data = 8'he3;
      17'd40843: data = 8'he0;
      17'd40844: data = 8'hde;
      17'd40845: data = 8'hdb;
      17'd40846: data = 8'hd8;
      17'd40847: data = 8'hd8;
      17'd40848: data = 8'hdb;
      17'd40849: data = 8'hd8;
      17'd40850: data = 8'hd3;
      17'd40851: data = 8'hd8;
      17'd40852: data = 8'hd8;
      17'd40853: data = 8'hd6;
      17'd40854: data = 8'hda;
      17'd40855: data = 8'hda;
      17'd40856: data = 8'he0;
      17'd40857: data = 8'he5;
      17'd40858: data = 8'heb;
      17'd40859: data = 8'hec;
      17'd40860: data = 8'hef;
      17'd40861: data = 8'hf5;
      17'd40862: data = 8'hfa;
      17'd40863: data = 8'hfe;
      17'd40864: data = 8'h01;
      17'd40865: data = 8'h05;
      17'd40866: data = 8'h05;
      17'd40867: data = 8'h0c;
      17'd40868: data = 8'h15;
      17'd40869: data = 8'h15;
      17'd40870: data = 8'h16;
      17'd40871: data = 8'h16;
      17'd40872: data = 8'h15;
      17'd40873: data = 8'h1b;
      17'd40874: data = 8'h22;
      17'd40875: data = 8'h22;
      17'd40876: data = 8'h1f;
      17'd40877: data = 8'h1f;
      17'd40878: data = 8'h1f;
      17'd40879: data = 8'h22;
      17'd40880: data = 8'h1f;
      17'd40881: data = 8'h19;
      17'd40882: data = 8'h13;
      17'd40883: data = 8'h13;
      17'd40884: data = 8'h15;
      17'd40885: data = 8'h12;
      17'd40886: data = 8'h05;
      17'd40887: data = 8'h04;
      17'd40888: data = 8'h02;
      17'd40889: data = 8'h00;
      17'd40890: data = 8'hfd;
      17'd40891: data = 8'hf6;
      17'd40892: data = 8'hf1;
      17'd40893: data = 8'hef;
      17'd40894: data = 8'hef;
      17'd40895: data = 8'hf1;
      17'd40896: data = 8'heb;
      17'd40897: data = 8'he4;
      17'd40898: data = 8'he4;
      17'd40899: data = 8'he3;
      17'd40900: data = 8'he3;
      17'd40901: data = 8'he3;
      17'd40902: data = 8'he4;
      17'd40903: data = 8'hde;
      17'd40904: data = 8'he3;
      17'd40905: data = 8'heb;
      17'd40906: data = 8'he5;
      17'd40907: data = 8'he9;
      17'd40908: data = 8'he7;
      17'd40909: data = 8'hec;
      17'd40910: data = 8'hf5;
      17'd40911: data = 8'hf5;
      17'd40912: data = 8'hf5;
      17'd40913: data = 8'hfd;
      17'd40914: data = 8'h02;
      17'd40915: data = 8'h04;
      17'd40916: data = 8'h09;
      17'd40917: data = 8'h05;
      17'd40918: data = 8'h06;
      17'd40919: data = 8'h0a;
      17'd40920: data = 8'h11;
      17'd40921: data = 8'h11;
      17'd40922: data = 8'h0c;
      17'd40923: data = 8'h0c;
      17'd40924: data = 8'h12;
      17'd40925: data = 8'h12;
      17'd40926: data = 8'h11;
      17'd40927: data = 8'h0a;
      17'd40928: data = 8'h06;
      17'd40929: data = 8'h0a;
      17'd40930: data = 8'h0c;
      17'd40931: data = 8'h0a;
      17'd40932: data = 8'h04;
      17'd40933: data = 8'h00;
      17'd40934: data = 8'hfe;
      17'd40935: data = 8'h00;
      17'd40936: data = 8'hf9;
      17'd40937: data = 8'hf6;
      17'd40938: data = 8'hf5;
      17'd40939: data = 8'hef;
      17'd40940: data = 8'hed;
      17'd40941: data = 8'hed;
      17'd40942: data = 8'hed;
      17'd40943: data = 8'he9;
      17'd40944: data = 8'heb;
      17'd40945: data = 8'hec;
      17'd40946: data = 8'he4;
      17'd40947: data = 8'hdb;
      17'd40948: data = 8'he0;
      17'd40949: data = 8'hd6;
      17'd40950: data = 8'hd5;
      17'd40951: data = 8'he5;
      17'd40952: data = 8'heb;
      17'd40953: data = 8'he9;
      17'd40954: data = 8'he9;
      17'd40955: data = 8'hf2;
      17'd40956: data = 8'hef;
      17'd40957: data = 8'hf4;
      17'd40958: data = 8'h02;
      17'd40959: data = 8'hfe;
      17'd40960: data = 8'hfc;
      17'd40961: data = 8'h04;
      17'd40962: data = 8'h06;
      17'd40963: data = 8'h00;
      17'd40964: data = 8'h04;
      17'd40965: data = 8'h09;
      17'd40966: data = 8'h00;
      17'd40967: data = 8'hfe;
      17'd40968: data = 8'h0c;
      17'd40969: data = 8'h0a;
      17'd40970: data = 8'h06;
      17'd40971: data = 8'h13;
      17'd40972: data = 8'h1b;
      17'd40973: data = 8'h13;
      17'd40974: data = 8'h0e;
      17'd40975: data = 8'h0d;
      17'd40976: data = 8'h09;
      17'd40977: data = 8'h05;
      17'd40978: data = 8'h0a;
      17'd40979: data = 8'h0a;
      17'd40980: data = 8'h01;
      17'd40981: data = 8'h00;
      17'd40982: data = 8'h04;
      17'd40983: data = 8'hfd;
      17'd40984: data = 8'hfa;
      17'd40985: data = 8'hfd;
      17'd40986: data = 8'hfa;
      17'd40987: data = 8'hf9;
      17'd40988: data = 8'h01;
      17'd40989: data = 8'h01;
      17'd40990: data = 8'hf9;
      17'd40991: data = 8'hfd;
      17'd40992: data = 8'hfd;
      17'd40993: data = 8'hf9;
      17'd40994: data = 8'hf4;
      17'd40995: data = 8'hf2;
      17'd40996: data = 8'hef;
      17'd40997: data = 8'hf4;
      17'd40998: data = 8'hfe;
      17'd40999: data = 8'hfe;
      17'd41000: data = 8'hf4;
      17'd41001: data = 8'hf4;
      17'd41002: data = 8'hfc;
      17'd41003: data = 8'hfc;
      17'd41004: data = 8'h00;
      17'd41005: data = 8'h01;
      17'd41006: data = 8'hfa;
      17'd41007: data = 8'h02;
      17'd41008: data = 8'h09;
      17'd41009: data = 8'h04;
      17'd41010: data = 8'h01;
      17'd41011: data = 8'h01;
      17'd41012: data = 8'h04;
      17'd41013: data = 8'h05;
      17'd41014: data = 8'h06;
      17'd41015: data = 8'h0c;
      17'd41016: data = 8'h0c;
      17'd41017: data = 8'h12;
      17'd41018: data = 8'h13;
      17'd41019: data = 8'h12;
      17'd41020: data = 8'h11;
      17'd41021: data = 8'h13;
      17'd41022: data = 8'h12;
      17'd41023: data = 8'h0d;
      17'd41024: data = 8'h13;
      17'd41025: data = 8'h15;
      17'd41026: data = 8'h0d;
      17'd41027: data = 8'h09;
      17'd41028: data = 8'h05;
      17'd41029: data = 8'h09;
      17'd41030: data = 8'h09;
      17'd41031: data = 8'h04;
      17'd41032: data = 8'h09;
      17'd41033: data = 8'hfe;
      17'd41034: data = 8'h06;
      17'd41035: data = 8'h0e;
      17'd41036: data = 8'h09;
      17'd41037: data = 8'h06;
      17'd41038: data = 8'h05;
      17'd41039: data = 8'h09;
      17'd41040: data = 8'h01;
      17'd41041: data = 8'h0a;
      17'd41042: data = 8'h02;
      17'd41043: data = 8'h01;
      17'd41044: data = 8'h06;
      17'd41045: data = 8'h04;
      17'd41046: data = 8'h0a;
      17'd41047: data = 8'h0c;
      17'd41048: data = 8'h0e;
      17'd41049: data = 8'h0a;
      17'd41050: data = 8'h0c;
      17'd41051: data = 8'h0e;
      17'd41052: data = 8'h12;
      17'd41053: data = 8'h0a;
      17'd41054: data = 8'h11;
      17'd41055: data = 8'h11;
      17'd41056: data = 8'h09;
      17'd41057: data = 8'h11;
      17'd41058: data = 8'h0d;
      17'd41059: data = 8'h0e;
      17'd41060: data = 8'h0c;
      17'd41061: data = 8'h13;
      17'd41062: data = 8'h13;
      17'd41063: data = 8'h06;
      17'd41064: data = 8'h02;
      17'd41065: data = 8'h09;
      17'd41066: data = 8'h01;
      17'd41067: data = 8'h01;
      17'd41068: data = 8'h06;
      17'd41069: data = 8'hfd;
      17'd41070: data = 8'hfe;
      17'd41071: data = 8'hfd;
      17'd41072: data = 8'h00;
      17'd41073: data = 8'hf4;
      17'd41074: data = 8'hfc;
      17'd41075: data = 8'h02;
      17'd41076: data = 8'hf9;
      17'd41077: data = 8'hfd;
      17'd41078: data = 8'hfc;
      17'd41079: data = 8'hfd;
      17'd41080: data = 8'h00;
      17'd41081: data = 8'h05;
      17'd41082: data = 8'h0d;
      17'd41083: data = 8'hfe;
      17'd41084: data = 8'hfa;
      17'd41085: data = 8'h05;
      17'd41086: data = 8'h02;
      17'd41087: data = 8'h06;
      17'd41088: data = 8'h05;
      17'd41089: data = 8'h06;
      17'd41090: data = 8'h01;
      17'd41091: data = 8'h05;
      17'd41092: data = 8'h0a;
      17'd41093: data = 8'hfe;
      17'd41094: data = 8'hfe;
      17'd41095: data = 8'h05;
      17'd41096: data = 8'h05;
      17'd41097: data = 8'hfd;
      17'd41098: data = 8'hfe;
      17'd41099: data = 8'hfd;
      17'd41100: data = 8'hfc;
      17'd41101: data = 8'hfa;
      17'd41102: data = 8'hfc;
      17'd41103: data = 8'hf2;
      17'd41104: data = 8'he9;
      17'd41105: data = 8'hed;
      17'd41106: data = 8'hec;
      17'd41107: data = 8'hed;
      17'd41108: data = 8'hec;
      17'd41109: data = 8'he7;
      17'd41110: data = 8'he4;
      17'd41111: data = 8'hdc;
      17'd41112: data = 8'hde;
      17'd41113: data = 8'he2;
      17'd41114: data = 8'hde;
      17'd41115: data = 8'he4;
      17'd41116: data = 8'he2;
      17'd41117: data = 8'he2;
      17'd41118: data = 8'he5;
      17'd41119: data = 8'he5;
      17'd41120: data = 8'he5;
      17'd41121: data = 8'he5;
      17'd41122: data = 8'hec;
      17'd41123: data = 8'heb;
      17'd41124: data = 8'hf1;
      17'd41125: data = 8'hf9;
      17'd41126: data = 8'hf4;
      17'd41127: data = 8'hf6;
      17'd41128: data = 8'h00;
      17'd41129: data = 8'h04;
      17'd41130: data = 8'hfe;
      17'd41131: data = 8'h02;
      17'd41132: data = 8'h0a;
      17'd41133: data = 8'h09;
      17'd41134: data = 8'h0d;
      17'd41135: data = 8'h13;
      17'd41136: data = 8'h12;
      17'd41137: data = 8'h12;
      17'd41138: data = 8'h12;
      17'd41139: data = 8'h12;
      17'd41140: data = 8'h12;
      17'd41141: data = 8'h13;
      17'd41142: data = 8'h15;
      17'd41143: data = 8'h15;
      17'd41144: data = 8'h12;
      17'd41145: data = 8'h11;
      17'd41146: data = 8'h13;
      17'd41147: data = 8'h11;
      17'd41148: data = 8'h0d;
      17'd41149: data = 8'h0a;
      17'd41150: data = 8'h06;
      17'd41151: data = 8'h05;
      17'd41152: data = 8'h09;
      17'd41153: data = 8'h01;
      17'd41154: data = 8'hfe;
      17'd41155: data = 8'hfe;
      17'd41156: data = 8'hfa;
      17'd41157: data = 8'hf9;
      17'd41158: data = 8'hf6;
      17'd41159: data = 8'hf4;
      17'd41160: data = 8'hef;
      17'd41161: data = 8'hf1;
      17'd41162: data = 8'hf4;
      17'd41163: data = 8'hf2;
      17'd41164: data = 8'hef;
      17'd41165: data = 8'hf1;
      17'd41166: data = 8'hf2;
      17'd41167: data = 8'hf1;
      17'd41168: data = 8'hf1;
      17'd41169: data = 8'hf2;
      17'd41170: data = 8'hf4;
      17'd41171: data = 8'hf4;
      17'd41172: data = 8'hf9;
      17'd41173: data = 8'hf6;
      17'd41174: data = 8'hfa;
      17'd41175: data = 8'hfc;
      17'd41176: data = 8'hfd;
      17'd41177: data = 8'h00;
      17'd41178: data = 8'h01;
      17'd41179: data = 8'h04;
      17'd41180: data = 8'h06;
      17'd41181: data = 8'h06;
      17'd41182: data = 8'h09;
      17'd41183: data = 8'h09;
      17'd41184: data = 8'h0a;
      17'd41185: data = 8'h0e;
      17'd41186: data = 8'h0a;
      17'd41187: data = 8'h04;
      17'd41188: data = 8'h05;
      17'd41189: data = 8'h0d;
      17'd41190: data = 8'h0a;
      17'd41191: data = 8'h06;
      17'd41192: data = 8'h06;
      17'd41193: data = 8'h01;
      17'd41194: data = 8'h01;
      17'd41195: data = 8'h04;
      17'd41196: data = 8'h02;
      17'd41197: data = 8'hfc;
      17'd41198: data = 8'hfa;
      17'd41199: data = 8'hf6;
      17'd41200: data = 8'hfa;
      17'd41201: data = 8'hfa;
      17'd41202: data = 8'hf4;
      17'd41203: data = 8'hf1;
      17'd41204: data = 8'hef;
      17'd41205: data = 8'hef;
      17'd41206: data = 8'hf1;
      17'd41207: data = 8'hed;
      17'd41208: data = 8'heb;
      17'd41209: data = 8'hed;
      17'd41210: data = 8'hed;
      17'd41211: data = 8'hf4;
      17'd41212: data = 8'hf6;
      17'd41213: data = 8'hf4;
      17'd41214: data = 8'he7;
      17'd41215: data = 8'he3;
      17'd41216: data = 8'he9;
      17'd41217: data = 8'he4;
      17'd41218: data = 8'heb;
      17'd41219: data = 8'hf5;
      17'd41220: data = 8'hf6;
      17'd41221: data = 8'hf1;
      17'd41222: data = 8'hf9;
      17'd41223: data = 8'h01;
      17'd41224: data = 8'h02;
      17'd41225: data = 8'h0a;
      17'd41226: data = 8'h09;
      17'd41227: data = 8'h06;
      17'd41228: data = 8'h06;
      17'd41229: data = 8'h0e;
      17'd41230: data = 8'h11;
      17'd41231: data = 8'h0a;
      17'd41232: data = 8'h01;
      17'd41233: data = 8'h05;
      17'd41234: data = 8'h09;
      17'd41235: data = 8'hf9;
      17'd41236: data = 8'hfe;
      17'd41237: data = 8'h06;
      17'd41238: data = 8'h04;
      17'd41239: data = 8'h05;
      17'd41240: data = 8'h0e;
      17'd41241: data = 8'h05;
      17'd41242: data = 8'hfe;
      17'd41243: data = 8'h01;
      17'd41244: data = 8'h02;
      17'd41245: data = 8'hfd;
      17'd41246: data = 8'hf9;
      17'd41247: data = 8'hfd;
      17'd41248: data = 8'hf4;
      17'd41249: data = 8'hf2;
      17'd41250: data = 8'hf9;
      17'd41251: data = 8'hf2;
      17'd41252: data = 8'hec;
      17'd41253: data = 8'hef;
      17'd41254: data = 8'hf6;
      17'd41255: data = 8'hf1;
      17'd41256: data = 8'hf5;
      17'd41257: data = 8'hfd;
      17'd41258: data = 8'hfd;
      17'd41259: data = 8'hfc;
      17'd41260: data = 8'hfc;
      17'd41261: data = 8'hfd;
      17'd41262: data = 8'hf5;
      17'd41263: data = 8'hf9;
      17'd41264: data = 8'hfa;
      17'd41265: data = 8'hf9;
      17'd41266: data = 8'hfa;
      17'd41267: data = 8'hfc;
      17'd41268: data = 8'hfe;
      17'd41269: data = 8'hfd;
      17'd41270: data = 8'hfe;
      17'd41271: data = 8'h01;
      17'd41272: data = 8'h05;
      17'd41273: data = 8'h05;
      17'd41274: data = 8'h05;
      17'd41275: data = 8'h05;
      17'd41276: data = 8'h0c;
      17'd41277: data = 8'h12;
      17'd41278: data = 8'h0d;
      17'd41279: data = 8'h06;
      17'd41280: data = 8'h06;
      17'd41281: data = 8'h06;
      17'd41282: data = 8'h0a;
      17'd41283: data = 8'h0e;
      17'd41284: data = 8'h09;
      17'd41285: data = 8'h05;
      17'd41286: data = 8'h0a;
      17'd41287: data = 8'h13;
      17'd41288: data = 8'h11;
      17'd41289: data = 8'h0e;
      17'd41290: data = 8'h0c;
      17'd41291: data = 8'h09;
      17'd41292: data = 8'h12;
      17'd41293: data = 8'h12;
      17'd41294: data = 8'h16;
      17'd41295: data = 8'h05;
      17'd41296: data = 8'h0c;
      17'd41297: data = 8'h13;
      17'd41298: data = 8'h09;
      17'd41299: data = 8'h09;
      17'd41300: data = 8'h0a;
      17'd41301: data = 8'h06;
      17'd41302: data = 8'h02;
      17'd41303: data = 8'h15;
      17'd41304: data = 8'h11;
      17'd41305: data = 8'h06;
      17'd41306: data = 8'h0e;
      17'd41307: data = 8'h1a;
      17'd41308: data = 8'h0a;
      17'd41309: data = 8'h0e;
      17'd41310: data = 8'h15;
      17'd41311: data = 8'h0a;
      17'd41312: data = 8'h0d;
      17'd41313: data = 8'h11;
      17'd41314: data = 8'h1b;
      17'd41315: data = 8'h0a;
      17'd41316: data = 8'h0c;
      17'd41317: data = 8'h0d;
      17'd41318: data = 8'h13;
      17'd41319: data = 8'h0d;
      17'd41320: data = 8'h09;
      17'd41321: data = 8'h13;
      17'd41322: data = 8'hfe;
      17'd41323: data = 8'h09;
      17'd41324: data = 8'h15;
      17'd41325: data = 8'h0e;
      17'd41326: data = 8'hfd;
      17'd41327: data = 8'h01;
      17'd41328: data = 8'hfd;
      17'd41329: data = 8'hef;
      17'd41330: data = 8'hfc;
      17'd41331: data = 8'hfe;
      17'd41332: data = 8'hfc;
      17'd41333: data = 8'hfc;
      17'd41334: data = 8'h06;
      17'd41335: data = 8'h04;
      17'd41336: data = 8'h00;
      17'd41337: data = 8'hfa;
      17'd41338: data = 8'h01;
      17'd41339: data = 8'h00;
      17'd41340: data = 8'hfe;
      17'd41341: data = 8'h06;
      17'd41342: data = 8'h05;
      17'd41343: data = 8'hfc;
      17'd41344: data = 8'h02;
      17'd41345: data = 8'h11;
      17'd41346: data = 8'h02;
      17'd41347: data = 8'h01;
      17'd41348: data = 8'h01;
      17'd41349: data = 8'h04;
      17'd41350: data = 8'h06;
      17'd41351: data = 8'h13;
      17'd41352: data = 8'h12;
      17'd41353: data = 8'h0c;
      17'd41354: data = 8'h0c;
      17'd41355: data = 8'h0c;
      17'd41356: data = 8'h0d;
      17'd41357: data = 8'h05;
      17'd41358: data = 8'h00;
      17'd41359: data = 8'hfe;
      17'd41360: data = 8'h01;
      17'd41361: data = 8'h04;
      17'd41362: data = 8'h02;
      17'd41363: data = 8'hf6;
      17'd41364: data = 8'hf1;
      17'd41365: data = 8'hf2;
      17'd41366: data = 8'hf4;
      17'd41367: data = 8'hec;
      17'd41368: data = 8'he7;
      17'd41369: data = 8'hef;
      17'd41370: data = 8'he9;
      17'd41371: data = 8'hef;
      17'd41372: data = 8'heb;
      17'd41373: data = 8'he5;
      17'd41374: data = 8'he2;
      17'd41375: data = 8'hde;
      17'd41376: data = 8'he0;
      17'd41377: data = 8'hdc;
      17'd41378: data = 8'hd8;
      17'd41379: data = 8'hdb;
      17'd41380: data = 8'hde;
      17'd41381: data = 8'hdc;
      17'd41382: data = 8'he3;
      17'd41383: data = 8'he3;
      17'd41384: data = 8'he0;
      17'd41385: data = 8'he2;
      17'd41386: data = 8'he9;
      17'd41387: data = 8'hed;
      17'd41388: data = 8'hef;
      17'd41389: data = 8'hfa;
      17'd41390: data = 8'hfd;
      17'd41391: data = 8'hfe;
      17'd41392: data = 8'hfe;
      17'd41393: data = 8'h02;
      17'd41394: data = 8'h04;
      17'd41395: data = 8'h04;
      17'd41396: data = 8'h04;
      17'd41397: data = 8'h06;
      17'd41398: data = 8'h09;
      17'd41399: data = 8'h0c;
      17'd41400: data = 8'h0c;
      17'd41401: data = 8'h0d;
      17'd41402: data = 8'h12;
      17'd41403: data = 8'h0d;
      17'd41404: data = 8'h0c;
      17'd41405: data = 8'h0e;
      17'd41406: data = 8'h0e;
      17'd41407: data = 8'h0d;
      17'd41408: data = 8'h11;
      17'd41409: data = 8'h12;
      17'd41410: data = 8'h09;
      17'd41411: data = 8'h06;
      17'd41412: data = 8'h05;
      17'd41413: data = 8'h01;
      17'd41414: data = 8'h02;
      17'd41415: data = 8'hfc;
      17'd41416: data = 8'hf9;
      17'd41417: data = 8'hfc;
      17'd41418: data = 8'hf9;
      17'd41419: data = 8'hf9;
      17'd41420: data = 8'hf4;
      17'd41421: data = 8'hf2;
      17'd41422: data = 8'hf2;
      17'd41423: data = 8'hf4;
      17'd41424: data = 8'hf2;
      17'd41425: data = 8'hef;
      17'd41426: data = 8'hf1;
      17'd41427: data = 8'hf2;
      17'd41428: data = 8'hf4;
      17'd41429: data = 8'hf5;
      17'd41430: data = 8'hef;
      17'd41431: data = 8'hf1;
      17'd41432: data = 8'hf4;
      17'd41433: data = 8'hf2;
      17'd41434: data = 8'hf6;
      17'd41435: data = 8'hfa;
      17'd41436: data = 8'hf9;
      17'd41437: data = 8'hf6;
      17'd41438: data = 8'h01;
      17'd41439: data = 8'h04;
      17'd41440: data = 8'h01;
      17'd41441: data = 8'h01;
      17'd41442: data = 8'h02;
      17'd41443: data = 8'h04;
      17'd41444: data = 8'h09;
      17'd41445: data = 8'h09;
      17'd41446: data = 8'h06;
      17'd41447: data = 8'h09;
      17'd41448: data = 8'h0a;
      17'd41449: data = 8'h09;
      17'd41450: data = 8'h05;
      17'd41451: data = 8'h04;
      17'd41452: data = 8'h02;
      17'd41453: data = 8'h01;
      17'd41454: data = 8'h04;
      17'd41455: data = 8'hfe;
      17'd41456: data = 8'hfc;
      17'd41457: data = 8'h00;
      17'd41458: data = 8'hfd;
      17'd41459: data = 8'hf6;
      17'd41460: data = 8'hf9;
      17'd41461: data = 8'hf5;
      17'd41462: data = 8'hf1;
      17'd41463: data = 8'hf1;
      17'd41464: data = 8'hf2;
      17'd41465: data = 8'hf2;
      17'd41466: data = 8'hed;
      17'd41467: data = 8'hef;
      17'd41468: data = 8'hec;
      17'd41469: data = 8'heb;
      17'd41470: data = 8'hec;
      17'd41471: data = 8'heb;
      17'd41472: data = 8'heb;
      17'd41473: data = 8'hec;
      17'd41474: data = 8'hf1;
      17'd41475: data = 8'hef;
      17'd41476: data = 8'hef;
      17'd41477: data = 8'hf6;
      17'd41478: data = 8'hfc;
      17'd41479: data = 8'hfd;
      17'd41480: data = 8'hf6;
      17'd41481: data = 8'hf4;
      17'd41482: data = 8'hf4;
      17'd41483: data = 8'hed;
      17'd41484: data = 8'hf4;
      17'd41485: data = 8'hfe;
      17'd41486: data = 8'hfe;
      17'd41487: data = 8'hfe;
      17'd41488: data = 8'hfc;
      17'd41489: data = 8'h00;
      17'd41490: data = 8'h00;
      17'd41491: data = 8'h05;
      17'd41492: data = 8'h0c;
      17'd41493: data = 8'h09;
      17'd41494: data = 8'h05;
      17'd41495: data = 8'h05;
      17'd41496: data = 8'h0c;
      17'd41497: data = 8'h0a;
      17'd41498: data = 8'h05;
      17'd41499: data = 8'h04;
      17'd41500: data = 8'hfe;
      17'd41501: data = 8'hfa;
      17'd41502: data = 8'hfc;
      17'd41503: data = 8'hfc;
      17'd41504: data = 8'hf9;
      17'd41505: data = 8'hfe;
      17'd41506: data = 8'h01;
      17'd41507: data = 8'h01;
      17'd41508: data = 8'hfe;
      17'd41509: data = 8'hf9;
      17'd41510: data = 8'hfc;
      17'd41511: data = 8'hfc;
      17'd41512: data = 8'hfc;
      17'd41513: data = 8'hf9;
      17'd41514: data = 8'hf5;
      17'd41515: data = 8'hf9;
      17'd41516: data = 8'hfa;
      17'd41517: data = 8'hfa;
      17'd41518: data = 8'hf5;
      17'd41519: data = 8'hf4;
      17'd41520: data = 8'hf6;
      17'd41521: data = 8'hfa;
      17'd41522: data = 8'hfc;
      17'd41523: data = 8'hfd;
      17'd41524: data = 8'h01;
      17'd41525: data = 8'h05;
      17'd41526: data = 8'h05;
      17'd41527: data = 8'h04;
      17'd41528: data = 8'h01;
      17'd41529: data = 8'h01;
      17'd41530: data = 8'h04;
      17'd41531: data = 8'h05;
      17'd41532: data = 8'h04;
      17'd41533: data = 8'h05;
      17'd41534: data = 8'h04;
      17'd41535: data = 8'h05;
      17'd41536: data = 8'h09;
      17'd41537: data = 8'h09;
      17'd41538: data = 8'h0a;
      17'd41539: data = 8'h09;
      17'd41540: data = 8'h0a;
      17'd41541: data = 8'h0a;
      17'd41542: data = 8'h0d;
      17'd41543: data = 8'h12;
      17'd41544: data = 8'h11;
      17'd41545: data = 8'h0d;
      17'd41546: data = 8'h09;
      17'd41547: data = 8'h0c;
      17'd41548: data = 8'h0c;
      17'd41549: data = 8'h0d;
      17'd41550: data = 8'h0c;
      17'd41551: data = 8'h0c;
      17'd41552: data = 8'h0c;
      17'd41553: data = 8'h0a;
      17'd41554: data = 8'h11;
      17'd41555: data = 8'h0c;
      17'd41556: data = 8'h0c;
      17'd41557: data = 8'h0c;
      17'd41558: data = 8'h09;
      17'd41559: data = 8'h11;
      17'd41560: data = 8'h0d;
      17'd41561: data = 8'h0d;
      17'd41562: data = 8'h11;
      17'd41563: data = 8'h11;
      17'd41564: data = 8'h09;
      17'd41565: data = 8'h0d;
      17'd41566: data = 8'h0a;
      17'd41567: data = 8'h09;
      17'd41568: data = 8'h0d;
      17'd41569: data = 8'h04;
      17'd41570: data = 8'h0e;
      17'd41571: data = 8'h0d;
      17'd41572: data = 8'h13;
      17'd41573: data = 8'h0e;
      17'd41574: data = 8'h0a;
      17'd41575: data = 8'h11;
      17'd41576: data = 8'h06;
      17'd41577: data = 8'h11;
      17'd41578: data = 8'h15;
      17'd41579: data = 8'h0d;
      17'd41580: data = 8'h13;
      17'd41581: data = 8'h13;
      17'd41582: data = 8'h06;
      17'd41583: data = 8'h0e;
      17'd41584: data = 8'h06;
      17'd41585: data = 8'h04;
      17'd41586: data = 8'h0c;
      17'd41587: data = 8'h0c;
      17'd41588: data = 8'h0d;
      17'd41589: data = 8'h06;
      17'd41590: data = 8'h11;
      17'd41591: data = 8'h02;
      17'd41592: data = 8'h06;
      17'd41593: data = 8'h06;
      17'd41594: data = 8'hfc;
      17'd41595: data = 8'h09;
      17'd41596: data = 8'h02;
      17'd41597: data = 8'h0a;
      17'd41598: data = 8'h04;
      17'd41599: data = 8'h06;
      17'd41600: data = 8'h04;
      17'd41601: data = 8'hfd;
      17'd41602: data = 8'h04;
      17'd41603: data = 8'h02;
      17'd41604: data = 8'h02;
      17'd41605: data = 8'hfd;
      17'd41606: data = 8'he7;
      17'd41607: data = 8'he0;
      17'd41608: data = 8'he4;
      17'd41609: data = 8'he5;
      17'd41610: data = 8'h02;
      17'd41611: data = 8'h05;
      17'd41612: data = 8'h06;
      17'd41613: data = 8'h0e;
      17'd41614: data = 8'h15;
      17'd41615: data = 8'h19;
      17'd41616: data = 8'h11;
      17'd41617: data = 8'h16;
      17'd41618: data = 8'h16;
      17'd41619: data = 8'h0a;
      17'd41620: data = 8'h0c;
      17'd41621: data = 8'h01;
      17'd41622: data = 8'hfa;
      17'd41623: data = 8'h05;
      17'd41624: data = 8'hfd;
      17'd41625: data = 8'hf9;
      17'd41626: data = 8'hed;
      17'd41627: data = 8'hef;
      17'd41628: data = 8'hf6;
      17'd41629: data = 8'hfd;
      17'd41630: data = 8'h09;
      17'd41631: data = 8'h06;
      17'd41632: data = 8'h09;
      17'd41633: data = 8'h05;
      17'd41634: data = 8'hfe;
      17'd41635: data = 8'hf9;
      17'd41636: data = 8'hef;
      17'd41637: data = 8'he7;
      17'd41638: data = 8'hec;
      17'd41639: data = 8'he2;
      17'd41640: data = 8'hde;
      17'd41641: data = 8'hde;
      17'd41642: data = 8'hda;
      17'd41643: data = 8'hde;
      17'd41644: data = 8'hd5;
      17'd41645: data = 8'hd6;
      17'd41646: data = 8'hd5;
      17'd41647: data = 8'hd6;
      17'd41648: data = 8'he4;
      17'd41649: data = 8'he7;
      17'd41650: data = 8'hf1;
      17'd41651: data = 8'hf4;
      17'd41652: data = 8'hec;
      17'd41653: data = 8'hec;
      17'd41654: data = 8'he9;
      17'd41655: data = 8'he7;
      17'd41656: data = 8'heb;
      17'd41657: data = 8'heb;
      17'd41658: data = 8'hf1;
      17'd41659: data = 8'hef;
      17'd41660: data = 8'hef;
      17'd41661: data = 8'hf6;
      17'd41662: data = 8'hf9;
      17'd41663: data = 8'hfe;
      17'd41664: data = 8'hfe;
      17'd41665: data = 8'hfd;
      17'd41666: data = 8'h05;
      17'd41667: data = 8'h0a;
      17'd41668: data = 8'h13;
      17'd41669: data = 8'h12;
      17'd41670: data = 8'h15;
      17'd41671: data = 8'h15;
      17'd41672: data = 8'h0c;
      17'd41673: data = 8'h0a;
      17'd41674: data = 8'h02;
      17'd41675: data = 8'h04;
      17'd41676: data = 8'h02;
      17'd41677: data = 8'h00;
      17'd41678: data = 8'h00;
      17'd41679: data = 8'hfa;
      17'd41680: data = 8'hfc;
      17'd41681: data = 8'hfd;
      17'd41682: data = 8'hfd;
      17'd41683: data = 8'hfd;
      17'd41684: data = 8'hf9;
      17'd41685: data = 8'hfa;
      17'd41686: data = 8'hfe;
      17'd41687: data = 8'hfe;
      17'd41688: data = 8'h02;
      17'd41689: data = 8'hfe;
      17'd41690: data = 8'hf5;
      17'd41691: data = 8'hf9;
      17'd41692: data = 8'hf4;
      17'd41693: data = 8'hef;
      17'd41694: data = 8'hec;
      17'd41695: data = 8'hec;
      17'd41696: data = 8'hed;
      17'd41697: data = 8'hf1;
      17'd41698: data = 8'hf4;
      17'd41699: data = 8'hf5;
      17'd41700: data = 8'hf6;
      17'd41701: data = 8'hfa;
      17'd41702: data = 8'hfe;
      17'd41703: data = 8'h01;
      17'd41704: data = 8'h02;
      17'd41705: data = 8'h04;
      17'd41706: data = 8'h0a;
      17'd41707: data = 8'h0c;
      17'd41708: data = 8'h0a;
      17'd41709: data = 8'h06;
      17'd41710: data = 8'h06;
      17'd41711: data = 8'h05;
      17'd41712: data = 8'h04;
      17'd41713: data = 8'h04;
      17'd41714: data = 8'h04;
      17'd41715: data = 8'h04;
      17'd41716: data = 8'h09;
      17'd41717: data = 8'h0a;
      17'd41718: data = 8'h09;
      17'd41719: data = 8'h0a;
      17'd41720: data = 8'h06;
      17'd41721: data = 8'h05;
      17'd41722: data = 8'h04;
      17'd41723: data = 8'h05;
      17'd41724: data = 8'h01;
      17'd41725: data = 8'h00;
      17'd41726: data = 8'h04;
      17'd41727: data = 8'hfc;
      17'd41728: data = 8'hf9;
      17'd41729: data = 8'hf6;
      17'd41730: data = 8'hf4;
      17'd41731: data = 8'hed;
      17'd41732: data = 8'hec;
      17'd41733: data = 8'hed;
      17'd41734: data = 8'hed;
      17'd41735: data = 8'hed;
      17'd41736: data = 8'hef;
      17'd41737: data = 8'hf1;
      17'd41738: data = 8'hed;
      17'd41739: data = 8'hf1;
      17'd41740: data = 8'hf1;
      17'd41741: data = 8'hf2;
      17'd41742: data = 8'hf4;
      17'd41743: data = 8'hf6;
      17'd41744: data = 8'hfa;
      17'd41745: data = 8'hf6;
      17'd41746: data = 8'hfa;
      17'd41747: data = 8'hfc;
      17'd41748: data = 8'hfc;
      17'd41749: data = 8'hfd;
      17'd41750: data = 8'hfa;
      17'd41751: data = 8'hf4;
      17'd41752: data = 8'hf4;
      17'd41753: data = 8'hf9;
      17'd41754: data = 8'hfd;
      17'd41755: data = 8'hfd;
      17'd41756: data = 8'hfa;
      17'd41757: data = 8'hfd;
      17'd41758: data = 8'h00;
      17'd41759: data = 8'h04;
      17'd41760: data = 8'h05;
      17'd41761: data = 8'h06;
      17'd41762: data = 8'h05;
      17'd41763: data = 8'h05;
      17'd41764: data = 8'h09;
      17'd41765: data = 8'h06;
      17'd41766: data = 8'h06;
      17'd41767: data = 8'h05;
      17'd41768: data = 8'h02;
      17'd41769: data = 8'h01;
      17'd41770: data = 8'hf6;
      17'd41771: data = 8'hf4;
      17'd41772: data = 8'hf6;
      17'd41773: data = 8'hf6;
      17'd41774: data = 8'hfc;
      17'd41775: data = 8'h00;
      17'd41776: data = 8'h00;
      17'd41777: data = 8'h00;
      17'd41778: data = 8'h04;
      17'd41779: data = 8'h05;
      17'd41780: data = 8'h04;
      17'd41781: data = 8'h05;
      17'd41782: data = 8'h05;
      17'd41783: data = 8'h04;
      17'd41784: data = 8'h04;
      17'd41785: data = 8'h01;
      17'd41786: data = 8'hfd;
      17'd41787: data = 8'hfd;
      17'd41788: data = 8'hf6;
      17'd41789: data = 8'hf6;
      17'd41790: data = 8'hf5;
      17'd41791: data = 8'hf5;
      17'd41792: data = 8'hfc;
      17'd41793: data = 8'hfd;
      17'd41794: data = 8'h01;
      17'd41795: data = 8'h05;
      17'd41796: data = 8'h09;
      17'd41797: data = 8'h04;
      17'd41798: data = 8'h01;
      17'd41799: data = 8'h05;
      17'd41800: data = 8'h04;
      17'd41801: data = 8'h05;
      17'd41802: data = 8'h04;
      17'd41803: data = 8'h02;
      17'd41804: data = 8'hfe;
      17'd41805: data = 8'h01;
      17'd41806: data = 8'h04;
      17'd41807: data = 8'h04;
      17'd41808: data = 8'h01;
      17'd41809: data = 8'h02;
      17'd41810: data = 8'h05;
      17'd41811: data = 8'h06;
      17'd41812: data = 8'h0c;
      17'd41813: data = 8'h0d;
      17'd41814: data = 8'h0d;
      17'd41815: data = 8'h0c;
      17'd41816: data = 8'h0d;
      17'd41817: data = 8'h0d;
      17'd41818: data = 8'h09;
      17'd41819: data = 8'h09;
      17'd41820: data = 8'h09;
      17'd41821: data = 8'h0a;
      17'd41822: data = 8'h0a;
      17'd41823: data = 8'h0c;
      17'd41824: data = 8'h0c;
      17'd41825: data = 8'h0c;
      17'd41826: data = 8'h0d;
      17'd41827: data = 8'h0e;
      17'd41828: data = 8'h0d;
      17'd41829: data = 8'h0d;
      17'd41830: data = 8'h0e;
      17'd41831: data = 8'h13;
      17'd41832: data = 8'h15;
      17'd41833: data = 8'h16;
      17'd41834: data = 8'h12;
      17'd41835: data = 8'h11;
      17'd41836: data = 8'h13;
      17'd41837: data = 8'h0d;
      17'd41838: data = 8'h0e;
      17'd41839: data = 8'h0d;
      17'd41840: data = 8'h0a;
      17'd41841: data = 8'h0a;
      17'd41842: data = 8'h0c;
      17'd41843: data = 8'h16;
      17'd41844: data = 8'h05;
      17'd41845: data = 8'h05;
      17'd41846: data = 8'h0e;
      17'd41847: data = 8'h05;
      17'd41848: data = 8'h04;
      17'd41849: data = 8'h11;
      17'd41850: data = 8'h09;
      17'd41851: data = 8'h01;
      17'd41852: data = 8'h12;
      17'd41853: data = 8'h0d;
      17'd41854: data = 8'h04;
      17'd41855: data = 8'h0a;
      17'd41856: data = 8'h09;
      17'd41857: data = 8'h02;
      17'd41858: data = 8'h0a;
      17'd41859: data = 8'h05;
      17'd41860: data = 8'h00;
      17'd41861: data = 8'h02;
      17'd41862: data = 8'h09;
      17'd41863: data = 8'h06;
      17'd41864: data = 8'hfc;
      17'd41865: data = 8'h05;
      17'd41866: data = 8'hfa;
      17'd41867: data = 8'h02;
      17'd41868: data = 8'h0c;
      17'd41869: data = 8'h01;
      17'd41870: data = 8'h0a;
      17'd41871: data = 8'h00;
      17'd41872: data = 8'h09;
      17'd41873: data = 8'h04;
      17'd41874: data = 8'h02;
      17'd41875: data = 8'h0a;
      17'd41876: data = 8'h00;
      17'd41877: data = 8'h05;
      17'd41878: data = 8'h0d;
      17'd41879: data = 8'hfd;
      17'd41880: data = 8'hf2;
      17'd41881: data = 8'hf4;
      17'd41882: data = 8'he3;
      17'd41883: data = 8'hf1;
      17'd41884: data = 8'hfa;
      17'd41885: data = 8'h02;
      17'd41886: data = 8'hfd;
      17'd41887: data = 8'h05;
      17'd41888: data = 8'h0d;
      17'd41889: data = 8'hf9;
      17'd41890: data = 8'h0e;
      17'd41891: data = 8'h05;
      17'd41892: data = 8'hf6;
      17'd41893: data = 8'hfd;
      17'd41894: data = 8'h09;
      17'd41895: data = 8'hf6;
      17'd41896: data = 8'hf4;
      17'd41897: data = 8'h01;
      17'd41898: data = 8'hf9;
      17'd41899: data = 8'heb;
      17'd41900: data = 8'hf1;
      17'd41901: data = 8'hf1;
      17'd41902: data = 8'he0;
      17'd41903: data = 8'hfa;
      17'd41904: data = 8'h01;
      17'd41905: data = 8'h04;
      17'd41906: data = 8'h02;
      17'd41907: data = 8'h09;
      17'd41908: data = 8'h05;
      17'd41909: data = 8'hf2;
      17'd41910: data = 8'hf5;
      17'd41911: data = 8'hf9;
      17'd41912: data = 8'hf4;
      17'd41913: data = 8'hf2;
      17'd41914: data = 8'hfd;
      17'd41915: data = 8'hf1;
      17'd41916: data = 8'hf1;
      17'd41917: data = 8'hef;
      17'd41918: data = 8'hf1;
      17'd41919: data = 8'heb;
      17'd41920: data = 8'he4;
      17'd41921: data = 8'hf1;
      17'd41922: data = 8'hf1;
      17'd41923: data = 8'hf4;
      17'd41924: data = 8'hf6;
      17'd41925: data = 8'hfd;
      17'd41926: data = 8'hfc;
      17'd41927: data = 8'hf6;
      17'd41928: data = 8'hf2;
      17'd41929: data = 8'hf2;
      17'd41930: data = 8'he3;
      17'd41931: data = 8'he9;
      17'd41932: data = 8'hf4;
      17'd41933: data = 8'hef;
      17'd41934: data = 8'hef;
      17'd41935: data = 8'hed;
      17'd41936: data = 8'hf4;
      17'd41937: data = 8'heb;
      17'd41938: data = 8'hf1;
      17'd41939: data = 8'hf4;
      17'd41940: data = 8'hef;
      17'd41941: data = 8'hf4;
      17'd41942: data = 8'hfe;
      17'd41943: data = 8'hfd;
      17'd41944: data = 8'hfc;
      17'd41945: data = 8'hfc;
      17'd41946: data = 8'hfe;
      17'd41947: data = 8'h00;
      17'd41948: data = 8'hf5;
      17'd41949: data = 8'hfa;
      17'd41950: data = 8'hf6;
      17'd41951: data = 8'hfa;
      17'd41952: data = 8'hfe;
      17'd41953: data = 8'h02;
      17'd41954: data = 8'h01;
      17'd41955: data = 8'hfe;
      17'd41956: data = 8'h01;
      17'd41957: data = 8'h01;
      17'd41958: data = 8'hfe;
      17'd41959: data = 8'h01;
      17'd41960: data = 8'h05;
      17'd41961: data = 8'h04;
      17'd41962: data = 8'h0a;
      17'd41963: data = 8'h09;
      17'd41964: data = 8'h09;
      17'd41965: data = 8'h04;
      17'd41966: data = 8'h06;
      17'd41967: data = 8'h04;
      17'd41968: data = 8'hfd;
      17'd41969: data = 8'hfe;
      17'd41970: data = 8'h01;
      17'd41971: data = 8'h02;
      17'd41972: data = 8'h02;
      17'd41973: data = 8'h04;
      17'd41974: data = 8'h00;
      17'd41975: data = 8'h00;
      17'd41976: data = 8'hfe;
      17'd41977: data = 8'hfe;
      17'd41978: data = 8'h00;
      17'd41979: data = 8'h00;
      17'd41980: data = 8'h01;
      17'd41981: data = 8'h00;
      17'd41982: data = 8'h04;
      17'd41983: data = 8'h01;
      17'd41984: data = 8'hfe;
      17'd41985: data = 8'hfd;
      17'd41986: data = 8'hfd;
      17'd41987: data = 8'hf9;
      17'd41988: data = 8'hf6;
      17'd41989: data = 8'hf9;
      17'd41990: data = 8'hf9;
      17'd41991: data = 8'hfd;
      17'd41992: data = 8'hfc;
      17'd41993: data = 8'hfa;
      17'd41994: data = 8'hfc;
      17'd41995: data = 8'hfa;
      17'd41996: data = 8'hfa;
      17'd41997: data = 8'hfd;
      17'd41998: data = 8'hfd;
      17'd41999: data = 8'hfd;
      17'd42000: data = 8'hfe;
      17'd42001: data = 8'h00;
      17'd42002: data = 8'h00;
      17'd42003: data = 8'hfe;
      17'd42004: data = 8'hfc;
      17'd42005: data = 8'hfa;
      17'd42006: data = 8'hfa;
      17'd42007: data = 8'hfc;
      17'd42008: data = 8'hfd;
      17'd42009: data = 8'hfd;
      17'd42010: data = 8'h00;
      17'd42011: data = 8'h01;
      17'd42012: data = 8'h00;
      17'd42013: data = 8'hfe;
      17'd42014: data = 8'h00;
      17'd42015: data = 8'h04;
      17'd42016: data = 8'h00;
      17'd42017: data = 8'hfc;
      17'd42018: data = 8'hfa;
      17'd42019: data = 8'hfd;
      17'd42020: data = 8'hfc;
      17'd42021: data = 8'hfe;
      17'd42022: data = 8'h01;
      17'd42023: data = 8'hf6;
      17'd42024: data = 8'hf2;
      17'd42025: data = 8'hf9;
      17'd42026: data = 8'hf6;
      17'd42027: data = 8'hf5;
      17'd42028: data = 8'hfd;
      17'd42029: data = 8'h01;
      17'd42030: data = 8'hf5;
      17'd42031: data = 8'hf6;
      17'd42032: data = 8'h00;
      17'd42033: data = 8'hfa;
      17'd42034: data = 8'hfa;
      17'd42035: data = 8'h02;
      17'd42036: data = 8'hfe;
      17'd42037: data = 8'hf2;
      17'd42038: data = 8'hfd;
      17'd42039: data = 8'h02;
      17'd42040: data = 8'hfc;
      17'd42041: data = 8'h00;
      17'd42042: data = 8'h04;
      17'd42043: data = 8'hfc;
      17'd42044: data = 8'hf6;
      17'd42045: data = 8'hfd;
      17'd42046: data = 8'hfe;
      17'd42047: data = 8'hfd;
      17'd42048: data = 8'h05;
      17'd42049: data = 8'h06;
      17'd42050: data = 8'hfe;
      17'd42051: data = 8'h00;
      17'd42052: data = 8'h01;
      17'd42053: data = 8'hfe;
      17'd42054: data = 8'h00;
      17'd42055: data = 8'h00;
      17'd42056: data = 8'hfe;
      17'd42057: data = 8'h00;
      17'd42058: data = 8'h01;
      17'd42059: data = 8'h00;
      17'd42060: data = 8'hfe;
      17'd42061: data = 8'hfe;
      17'd42062: data = 8'hfe;
      17'd42063: data = 8'hfc;
      17'd42064: data = 8'hfd;
      17'd42065: data = 8'hfc;
      17'd42066: data = 8'hfe;
      17'd42067: data = 8'h01;
      17'd42068: data = 8'h02;
      17'd42069: data = 8'h02;
      17'd42070: data = 8'h01;
      17'd42071: data = 8'h00;
      17'd42072: data = 8'h00;
      17'd42073: data = 8'h02;
      17'd42074: data = 8'h02;
      17'd42075: data = 8'h02;
      17'd42076: data = 8'h01;
      17'd42077: data = 8'h05;
      17'd42078: data = 8'h05;
      17'd42079: data = 8'h04;
      17'd42080: data = 8'h06;
      17'd42081: data = 8'h04;
      17'd42082: data = 8'h02;
      17'd42083: data = 8'h05;
      17'd42084: data = 8'h05;
      17'd42085: data = 8'h06;
      17'd42086: data = 8'h06;
      17'd42087: data = 8'h06;
      17'd42088: data = 8'h09;
      17'd42089: data = 8'h06;
      17'd42090: data = 8'h06;
      17'd42091: data = 8'h09;
      17'd42092: data = 8'h06;
      17'd42093: data = 8'h0a;
      17'd42094: data = 8'h0a;
      17'd42095: data = 8'h0c;
      17'd42096: data = 8'h0a;
      17'd42097: data = 8'h09;
      17'd42098: data = 8'h0c;
      17'd42099: data = 8'h0a;
      17'd42100: data = 8'h06;
      17'd42101: data = 8'h04;
      17'd42102: data = 8'h05;
      17'd42103: data = 8'h0a;
      17'd42104: data = 8'h0a;
      17'd42105: data = 8'h0a;
      17'd42106: data = 8'h09;
      17'd42107: data = 8'h0d;
      17'd42108: data = 8'h0c;
      17'd42109: data = 8'h0c;
      17'd42110: data = 8'h0a;
      17'd42111: data = 8'h0a;
      17'd42112: data = 8'h0e;
      17'd42113: data = 8'h0c;
      17'd42114: data = 8'h0a;
      17'd42115: data = 8'h11;
      17'd42116: data = 8'h0d;
      17'd42117: data = 8'h05;
      17'd42118: data = 8'h0a;
      17'd42119: data = 8'h06;
      17'd42120: data = 8'h01;
      17'd42121: data = 8'h01;
      17'd42122: data = 8'h0a;
      17'd42123: data = 8'h04;
      17'd42124: data = 8'h00;
      17'd42125: data = 8'h0d;
      17'd42126: data = 8'h05;
      17'd42127: data = 8'h04;
      17'd42128: data = 8'h13;
      17'd42129: data = 8'h02;
      17'd42130: data = 8'h04;
      17'd42131: data = 8'h06;
      17'd42132: data = 8'h04;
      17'd42133: data = 8'h0d;
      17'd42134: data = 8'hfe;
      17'd42135: data = 8'h06;
      17'd42136: data = 8'h06;
      17'd42137: data = 8'hf6;
      17'd42138: data = 8'h0c;
      17'd42139: data = 8'h06;
      17'd42140: data = 8'h00;
      17'd42141: data = 8'h0c;
      17'd42142: data = 8'hfe;
      17'd42143: data = 8'h06;
      17'd42144: data = 8'h04;
      17'd42145: data = 8'h04;
      17'd42146: data = 8'h0c;
      17'd42147: data = 8'hf2;
      17'd42148: data = 8'h09;
      17'd42149: data = 8'h02;
      17'd42150: data = 8'hf6;
      17'd42151: data = 8'h06;
      17'd42152: data = 8'hfa;
      17'd42153: data = 8'hf6;
      17'd42154: data = 8'h00;
      17'd42155: data = 8'hf9;
      17'd42156: data = 8'hfe;
      17'd42157: data = 8'hf6;
      17'd42158: data = 8'hf5;
      17'd42159: data = 8'h06;
      17'd42160: data = 8'hfa;
      17'd42161: data = 8'h01;
      17'd42162: data = 8'hfa;
      17'd42163: data = 8'hf5;
      17'd42164: data = 8'hfa;
      17'd42165: data = 8'hfc;
      17'd42166: data = 8'h01;
      17'd42167: data = 8'hf2;
      17'd42168: data = 8'hf6;
      17'd42169: data = 8'h00;
      17'd42170: data = 8'h01;
      17'd42171: data = 8'hfa;
      17'd42172: data = 8'hfd;
      17'd42173: data = 8'hf2;
      17'd42174: data = 8'hf4;
      17'd42175: data = 8'hf4;
      17'd42176: data = 8'hfd;
      17'd42177: data = 8'hfa;
      17'd42178: data = 8'hed;
      17'd42179: data = 8'h00;
      17'd42180: data = 8'hfa;
      17'd42181: data = 8'hf5;
      17'd42182: data = 8'hfa;
      17'd42183: data = 8'h00;
      17'd42184: data = 8'hf9;
      17'd42185: data = 8'hfc;
      17'd42186: data = 8'hfe;
      17'd42187: data = 8'h01;
      17'd42188: data = 8'hf6;
      17'd42189: data = 8'hfe;
      17'd42190: data = 8'h0a;
      17'd42191: data = 8'hf9;
      17'd42192: data = 8'hfe;
      17'd42193: data = 8'hfe;
      17'd42194: data = 8'hfd;
      17'd42195: data = 8'hf6;
      17'd42196: data = 8'hfd;
      17'd42197: data = 8'h02;
      17'd42198: data = 8'hfc;
      17'd42199: data = 8'hf9;
      17'd42200: data = 8'hfd;
      17'd42201: data = 8'hf5;
      17'd42202: data = 8'hf2;
      17'd42203: data = 8'hfd;
      17'd42204: data = 8'hf4;
      17'd42205: data = 8'hf5;
      17'd42206: data = 8'hf1;
      17'd42207: data = 8'hf5;
      17'd42208: data = 8'hf2;
      17'd42209: data = 8'hf1;
      17'd42210: data = 8'hf2;
      17'd42211: data = 8'hf1;
      17'd42212: data = 8'hec;
      17'd42213: data = 8'hed;
      17'd42214: data = 8'hef;
      17'd42215: data = 8'heb;
      17'd42216: data = 8'hef;
      17'd42217: data = 8'hec;
      17'd42218: data = 8'hf5;
      17'd42219: data = 8'hec;
      17'd42220: data = 8'hed;
      17'd42221: data = 8'hf1;
      17'd42222: data = 8'hed;
      17'd42223: data = 8'hf2;
      17'd42224: data = 8'hf2;
      17'd42225: data = 8'hf5;
      17'd42226: data = 8'hf4;
      17'd42227: data = 8'hf5;
      17'd42228: data = 8'hf5;
      17'd42229: data = 8'hf9;
      17'd42230: data = 8'hf4;
      17'd42231: data = 8'hfd;
      17'd42232: data = 8'hf9;
      17'd42233: data = 8'hf6;
      17'd42234: data = 8'hfd;
      17'd42235: data = 8'hfe;
      17'd42236: data = 8'h01;
      17'd42237: data = 8'hfe;
      17'd42238: data = 8'h01;
      17'd42239: data = 8'h01;
      17'd42240: data = 8'h02;
      17'd42241: data = 8'h01;
      17'd42242: data = 8'h01;
      17'd42243: data = 8'hfe;
      17'd42244: data = 8'h06;
      17'd42245: data = 8'h04;
      17'd42246: data = 8'h02;
      17'd42247: data = 8'h04;
      17'd42248: data = 8'h02;
      17'd42249: data = 8'h09;
      17'd42250: data = 8'h01;
      17'd42251: data = 8'h04;
      17'd42252: data = 8'h04;
      17'd42253: data = 8'h00;
      17'd42254: data = 8'h05;
      17'd42255: data = 8'h06;
      17'd42256: data = 8'h02;
      17'd42257: data = 8'h01;
      17'd42258: data = 8'h02;
      17'd42259: data = 8'h05;
      17'd42260: data = 8'h01;
      17'd42261: data = 8'h00;
      17'd42262: data = 8'h02;
      17'd42263: data = 8'hfe;
      17'd42264: data = 8'h04;
      17'd42265: data = 8'h01;
      17'd42266: data = 8'h00;
      17'd42267: data = 8'h00;
      17'd42268: data = 8'h00;
      17'd42269: data = 8'h02;
      17'd42270: data = 8'h02;
      17'd42271: data = 8'h01;
      17'd42272: data = 8'h01;
      17'd42273: data = 8'h01;
      17'd42274: data = 8'h01;
      17'd42275: data = 8'h04;
      17'd42276: data = 8'h05;
      17'd42277: data = 8'h05;
      17'd42278: data = 8'h01;
      17'd42279: data = 8'h02;
      17'd42280: data = 8'h00;
      17'd42281: data = 8'h01;
      17'd42282: data = 8'h02;
      17'd42283: data = 8'h01;
      17'd42284: data = 8'h02;
      17'd42285: data = 8'h02;
      17'd42286: data = 8'h00;
      17'd42287: data = 8'h00;
      17'd42288: data = 8'h01;
      17'd42289: data = 8'h01;
      17'd42290: data = 8'h02;
      17'd42291: data = 8'h02;
      17'd42292: data = 8'h04;
      17'd42293: data = 8'hfe;
      17'd42294: data = 8'hfe;
      17'd42295: data = 8'h00;
      17'd42296: data = 8'hfd;
      17'd42297: data = 8'hfe;
      17'd42298: data = 8'hfe;
      17'd42299: data = 8'hfe;
      17'd42300: data = 8'hfd;
      17'd42301: data = 8'hfc;
      17'd42302: data = 8'hfc;
      17'd42303: data = 8'hfd;
      17'd42304: data = 8'hfc;
      17'd42305: data = 8'hfd;
      17'd42306: data = 8'hfc;
      17'd42307: data = 8'hf9;
      17'd42308: data = 8'hf9;
      17'd42309: data = 8'hfe;
      17'd42310: data = 8'hfd;
      17'd42311: data = 8'hfa;
      17'd42312: data = 8'hfd;
      17'd42313: data = 8'hfd;
      17'd42314: data = 8'hfa;
      17'd42315: data = 8'hfa;
      17'd42316: data = 8'h01;
      17'd42317: data = 8'hfe;
      17'd42318: data = 8'hfd;
      17'd42319: data = 8'h00;
      17'd42320: data = 8'h04;
      17'd42321: data = 8'hfd;
      17'd42322: data = 8'hfd;
      17'd42323: data = 8'h01;
      17'd42324: data = 8'hfe;
      17'd42325: data = 8'hfe;
      17'd42326: data = 8'h00;
      17'd42327: data = 8'hfc;
      17'd42328: data = 8'hfa;
      17'd42329: data = 8'hfe;
      17'd42330: data = 8'h00;
      17'd42331: data = 8'hfd;
      17'd42332: data = 8'hfd;
      17'd42333: data = 8'hfe;
      17'd42334: data = 8'hfd;
      17'd42335: data = 8'hfe;
      17'd42336: data = 8'hfe;
      17'd42337: data = 8'hfc;
      17'd42338: data = 8'hf9;
      17'd42339: data = 8'hfd;
      17'd42340: data = 8'hfe;
      17'd42341: data = 8'hfa;
      17'd42342: data = 8'hfa;
      17'd42343: data = 8'hfc;
      17'd42344: data = 8'hfc;
      17'd42345: data = 8'hfc;
      17'd42346: data = 8'hfd;
      17'd42347: data = 8'hfd;
      17'd42348: data = 8'hfd;
      17'd42349: data = 8'hfe;
      17'd42350: data = 8'h01;
      17'd42351: data = 8'h01;
      17'd42352: data = 8'hfe;
      17'd42353: data = 8'h01;
      17'd42354: data = 8'h02;
      17'd42355: data = 8'h02;
      17'd42356: data = 8'h04;
      17'd42357: data = 8'h04;
      17'd42358: data = 8'h00;
      17'd42359: data = 8'h01;
      17'd42360: data = 8'h05;
      17'd42361: data = 8'h09;
      17'd42362: data = 8'h05;
      17'd42363: data = 8'h02;
      17'd42364: data = 8'h06;
      17'd42365: data = 8'h06;
      17'd42366: data = 8'h05;
      17'd42367: data = 8'h09;
      17'd42368: data = 8'h09;
      17'd42369: data = 8'h05;
      17'd42370: data = 8'h06;
      17'd42371: data = 8'h0a;
      17'd42372: data = 8'h09;
      17'd42373: data = 8'h09;
      17'd42374: data = 8'h06;
      17'd42375: data = 8'h06;
      17'd42376: data = 8'h09;
      17'd42377: data = 8'h06;
      17'd42378: data = 8'h06;
      17'd42379: data = 8'h06;
      17'd42380: data = 8'h09;
      17'd42381: data = 8'h0c;
      17'd42382: data = 8'h0a;
      17'd42383: data = 8'h04;
      17'd42384: data = 8'h06;
      17'd42385: data = 8'h06;
      17'd42386: data = 8'h09;
      17'd42387: data = 8'h05;
      17'd42388: data = 8'h06;
      17'd42389: data = 8'h06;
      17'd42390: data = 8'h05;
      17'd42391: data = 8'h06;
      17'd42392: data = 8'h0a;
      17'd42393: data = 8'h06;
      17'd42394: data = 8'h0a;
      17'd42395: data = 8'h09;
      17'd42396: data = 8'h06;
      17'd42397: data = 8'h0a;
      17'd42398: data = 8'h06;
      17'd42399: data = 8'h0a;
      17'd42400: data = 8'h09;
      17'd42401: data = 8'h09;
      17'd42402: data = 8'h05;
      17'd42403: data = 8'h02;
      17'd42404: data = 8'h05;
      17'd42405: data = 8'h05;
      17'd42406: data = 8'h09;
      17'd42407: data = 8'h06;
      17'd42408: data = 8'h04;
      17'd42409: data = 8'h0a;
      17'd42410: data = 8'h06;
      17'd42411: data = 8'h05;
      17'd42412: data = 8'h06;
      17'd42413: data = 8'h01;
      17'd42414: data = 8'h05;
      17'd42415: data = 8'h09;
      17'd42416: data = 8'h04;
      17'd42417: data = 8'h01;
      17'd42418: data = 8'h04;
      17'd42419: data = 8'h05;
      17'd42420: data = 8'h05;
      17'd42421: data = 8'h0a;
      17'd42422: data = 8'h05;
      17'd42423: data = 8'h01;
      17'd42424: data = 8'h00;
      17'd42425: data = 8'h05;
      17'd42426: data = 8'h06;
      17'd42427: data = 8'hfd;
      17'd42428: data = 8'hfe;
      17'd42429: data = 8'h01;
      17'd42430: data = 8'hfd;
      17'd42431: data = 8'h01;
      17'd42432: data = 8'h01;
      17'd42433: data = 8'hfe;
      17'd42434: data = 8'h01;
      17'd42435: data = 8'h01;
      17'd42436: data = 8'h09;
      17'd42437: data = 8'h02;
      17'd42438: data = 8'h01;
      17'd42439: data = 8'h04;
      17'd42440: data = 8'hfc;
      17'd42441: data = 8'hfe;
      17'd42442: data = 8'hfa;
      17'd42443: data = 8'hfc;
      17'd42444: data = 8'hfd;
      17'd42445: data = 8'hf4;
      17'd42446: data = 8'hfd;
      17'd42447: data = 8'h04;
      17'd42448: data = 8'hf5;
      17'd42449: data = 8'hfa;
      17'd42450: data = 8'h06;
      17'd42451: data = 8'h00;
      17'd42452: data = 8'hf1;
      17'd42453: data = 8'hfc;
      17'd42454: data = 8'h02;
      17'd42455: data = 8'hf9;
      17'd42456: data = 8'hfe;
      17'd42457: data = 8'h04;
      17'd42458: data = 8'hf5;
      17'd42459: data = 8'hf1;
      17'd42460: data = 8'hfd;
      17'd42461: data = 8'hfc;
      17'd42462: data = 8'hf6;
      17'd42463: data = 8'hfc;
      17'd42464: data = 8'hfe;
      17'd42465: data = 8'hfe;
      17'd42466: data = 8'hfc;
      17'd42467: data = 8'hfe;
      17'd42468: data = 8'hf6;
      17'd42469: data = 8'hf2;
      17'd42470: data = 8'hfc;
      17'd42471: data = 8'hfa;
      17'd42472: data = 8'hf6;
      17'd42473: data = 8'hf9;
      17'd42474: data = 8'hf2;
      17'd42475: data = 8'hf6;
      17'd42476: data = 8'hfd;
      17'd42477: data = 8'hf1;
      17'd42478: data = 8'hf2;
      17'd42479: data = 8'hfa;
      17'd42480: data = 8'hf9;
      17'd42481: data = 8'hfd;
      17'd42482: data = 8'h04;
      17'd42483: data = 8'hf9;
      17'd42484: data = 8'hf6;
      17'd42485: data = 8'h01;
      17'd42486: data = 8'hfc;
      17'd42487: data = 8'hf1;
      17'd42488: data = 8'hf5;
      17'd42489: data = 8'hf9;
      17'd42490: data = 8'hf2;
      17'd42491: data = 8'hf9;
      17'd42492: data = 8'h00;
      17'd42493: data = 8'hf5;
      17'd42494: data = 8'hf6;
      17'd42495: data = 8'h02;
      17'd42496: data = 8'hfa;
      17'd42497: data = 8'hf5;
      17'd42498: data = 8'h00;
      17'd42499: data = 8'h02;
      17'd42500: data = 8'hfc;
      17'd42501: data = 8'hfd;
      17'd42502: data = 8'hfd;
      17'd42503: data = 8'hf9;
      17'd42504: data = 8'hf6;
      17'd42505: data = 8'hfc;
      17'd42506: data = 8'hf5;
      17'd42507: data = 8'hef;
      17'd42508: data = 8'hfa;
      17'd42509: data = 8'hfd;
      17'd42510: data = 8'hfa;
      17'd42511: data = 8'hf4;
      17'd42512: data = 8'hf4;
      17'd42513: data = 8'hf5;
      17'd42514: data = 8'hfa;
      17'd42515: data = 8'hfa;
      17'd42516: data = 8'hf6;
      17'd42517: data = 8'hf2;
      17'd42518: data = 8'hf1;
      17'd42519: data = 8'hf9;
      17'd42520: data = 8'hfd;
      17'd42521: data = 8'hf4;
      17'd42522: data = 8'hf1;
      17'd42523: data = 8'hf6;
      17'd42524: data = 8'hf5;
      17'd42525: data = 8'hf9;
      17'd42526: data = 8'hf6;
      17'd42527: data = 8'hf9;
      17'd42528: data = 8'hf6;
      17'd42529: data = 8'hfd;
      17'd42530: data = 8'h01;
      17'd42531: data = 8'hf6;
      17'd42532: data = 8'hfa;
      17'd42533: data = 8'hfc;
      17'd42534: data = 8'hfa;
      17'd42535: data = 8'hfc;
      17'd42536: data = 8'hfc;
      17'd42537: data = 8'hfa;
      17'd42538: data = 8'hfc;
      17'd42539: data = 8'h00;
      17'd42540: data = 8'h00;
      17'd42541: data = 8'hfd;
      17'd42542: data = 8'hfc;
      17'd42543: data = 8'hfe;
      17'd42544: data = 8'hfe;
      17'd42545: data = 8'h02;
      17'd42546: data = 8'h01;
      17'd42547: data = 8'h00;
      17'd42548: data = 8'hfd;
      17'd42549: data = 8'h00;
      17'd42550: data = 8'h01;
      17'd42551: data = 8'h00;
      17'd42552: data = 8'h00;
      17'd42553: data = 8'h02;
      17'd42554: data = 8'h02;
      17'd42555: data = 8'h01;
      17'd42556: data = 8'h05;
      17'd42557: data = 8'h05;
      17'd42558: data = 8'h05;
      17'd42559: data = 8'h04;
      17'd42560: data = 8'h01;
      17'd42561: data = 8'h01;
      17'd42562: data = 8'h00;
      17'd42563: data = 8'hfd;
      17'd42564: data = 8'h00;
      17'd42565: data = 8'h04;
      17'd42566: data = 8'hfe;
      17'd42567: data = 8'h02;
      17'd42568: data = 8'h05;
      17'd42569: data = 8'h00;
      17'd42570: data = 8'h01;
      17'd42571: data = 8'h04;
      17'd42572: data = 8'h01;
      17'd42573: data = 8'h00;
      17'd42574: data = 8'h02;
      17'd42575: data = 8'h04;
      17'd42576: data = 8'h02;
      17'd42577: data = 8'h01;
      17'd42578: data = 8'h02;
      17'd42579: data = 8'hfe;
      17'd42580: data = 8'hfd;
      17'd42581: data = 8'h00;
      17'd42582: data = 8'h00;
      17'd42583: data = 8'hfe;
      17'd42584: data = 8'h04;
      17'd42585: data = 8'h02;
      17'd42586: data = 8'hf9;
      17'd42587: data = 8'h00;
      17'd42588: data = 8'h01;
      17'd42589: data = 8'hfd;
      17'd42590: data = 8'h00;
      17'd42591: data = 8'h02;
      17'd42592: data = 8'h00;
      17'd42593: data = 8'h02;
      17'd42594: data = 8'h04;
      17'd42595: data = 8'h04;
      17'd42596: data = 8'h01;
      17'd42597: data = 8'hfd;
      17'd42598: data = 8'h00;
      17'd42599: data = 8'hfd;
      17'd42600: data = 8'hfc;
      17'd42601: data = 8'h00;
      17'd42602: data = 8'hfd;
      17'd42603: data = 8'hfd;
      17'd42604: data = 8'h00;
      17'd42605: data = 8'h00;
      17'd42606: data = 8'hfd;
      17'd42607: data = 8'hfd;
      17'd42608: data = 8'hfe;
      17'd42609: data = 8'hfe;
      17'd42610: data = 8'h00;
      17'd42611: data = 8'h00;
      17'd42612: data = 8'hfe;
      17'd42613: data = 8'hfe;
      17'd42614: data = 8'h00;
      17'd42615: data = 8'hfc;
      17'd42616: data = 8'hfd;
      17'd42617: data = 8'hfe;
      17'd42618: data = 8'hfc;
      17'd42619: data = 8'hfe;
      17'd42620: data = 8'h02;
      17'd42621: data = 8'h01;
      17'd42622: data = 8'h02;
      17'd42623: data = 8'h04;
      17'd42624: data = 8'h01;
      17'd42625: data = 8'h01;
      17'd42626: data = 8'h02;
      17'd42627: data = 8'h04;
      17'd42628: data = 8'h02;
      17'd42629: data = 8'h01;
      17'd42630: data = 8'h00;
      17'd42631: data = 8'hfe;
      17'd42632: data = 8'h01;
      17'd42633: data = 8'h01;
      17'd42634: data = 8'h01;
      17'd42635: data = 8'h00;
      17'd42636: data = 8'h00;
      17'd42637: data = 8'h04;
      17'd42638: data = 8'h04;
      17'd42639: data = 8'h01;
      17'd42640: data = 8'h02;
      17'd42641: data = 8'h01;
      17'd42642: data = 8'hfe;
      17'd42643: data = 8'h01;
      17'd42644: data = 8'h00;
      17'd42645: data = 8'hfd;
      17'd42646: data = 8'hfd;
      17'd42647: data = 8'hfd;
      17'd42648: data = 8'hfe;
      17'd42649: data = 8'hfe;
      17'd42650: data = 8'hfe;
      17'd42651: data = 8'h00;
      17'd42652: data = 8'h00;
      17'd42653: data = 8'h00;
      17'd42654: data = 8'h04;
      17'd42655: data = 8'h05;
      17'd42656: data = 8'h04;
      17'd42657: data = 8'h05;
      17'd42658: data = 8'h02;
      17'd42659: data = 8'h02;
      17'd42660: data = 8'h09;
      17'd42661: data = 8'h09;
      17'd42662: data = 8'h05;
      17'd42663: data = 8'h02;
      17'd42664: data = 8'h05;
      17'd42665: data = 8'h0c;
      17'd42666: data = 8'h0c;
      17'd42667: data = 8'h05;
      17'd42668: data = 8'h04;
      17'd42669: data = 8'h05;
      17'd42670: data = 8'h09;
      17'd42671: data = 8'h0a;
      17'd42672: data = 8'h09;
      17'd42673: data = 8'h04;
      17'd42674: data = 8'h04;
      17'd42675: data = 8'h05;
      17'd42676: data = 8'h0c;
      17'd42677: data = 8'h06;
      17'd42678: data = 8'h00;
      17'd42679: data = 8'h05;
      17'd42680: data = 8'h06;
      17'd42681: data = 8'h09;
      17'd42682: data = 8'h09;
      17'd42683: data = 8'h04;
      17'd42684: data = 8'h05;
      17'd42685: data = 8'h06;
      17'd42686: data = 8'h09;
      17'd42687: data = 8'h06;
      17'd42688: data = 8'h04;
      17'd42689: data = 8'h09;
      17'd42690: data = 8'h06;
      17'd42691: data = 8'h0a;
      17'd42692: data = 8'h0d;
      17'd42693: data = 8'h05;
      17'd42694: data = 8'h06;
      17'd42695: data = 8'h09;
      17'd42696: data = 8'h04;
      17'd42697: data = 8'h05;
      17'd42698: data = 8'h05;
      17'd42699: data = 8'h04;
      17'd42700: data = 8'h01;
      17'd42701: data = 8'h01;
      17'd42702: data = 8'h02;
      17'd42703: data = 8'hfd;
      17'd42704: data = 8'h02;
      17'd42705: data = 8'h06;
      17'd42706: data = 8'hfa;
      17'd42707: data = 8'hfd;
      17'd42708: data = 8'h04;
      17'd42709: data = 8'h00;
      17'd42710: data = 8'h00;
      17'd42711: data = 8'h01;
      17'd42712: data = 8'h01;
      17'd42713: data = 8'h00;
      17'd42714: data = 8'h00;
      17'd42715: data = 8'h05;
      17'd42716: data = 8'h04;
      17'd42717: data = 8'hfd;
      17'd42718: data = 8'h00;
      17'd42719: data = 8'h04;
      17'd42720: data = 8'h02;
      17'd42721: data = 8'hfe;
      17'd42722: data = 8'h01;
      17'd42723: data = 8'hfe;
      17'd42724: data = 8'hfd;
      17'd42725: data = 8'hfd;
      17'd42726: data = 8'hfe;
      17'd42727: data = 8'hfd;
      17'd42728: data = 8'hf9;
      17'd42729: data = 8'hfd;
      17'd42730: data = 8'h02;
      17'd42731: data = 8'h00;
      17'd42732: data = 8'h00;
      17'd42733: data = 8'hfe;
      17'd42734: data = 8'hfa;
      17'd42735: data = 8'hfe;
      17'd42736: data = 8'h04;
      17'd42737: data = 8'h01;
      17'd42738: data = 8'hfd;
      17'd42739: data = 8'h01;
      17'd42740: data = 8'hfc;
      17'd42741: data = 8'hf9;
      17'd42742: data = 8'h04;
      17'd42743: data = 8'hfe;
      17'd42744: data = 8'hf5;
      17'd42745: data = 8'hfc;
      17'd42746: data = 8'hfa;
      17'd42747: data = 8'hfa;
      17'd42748: data = 8'hfd;
      17'd42749: data = 8'h01;
      17'd42750: data = 8'h01;
      17'd42751: data = 8'hf4;
      17'd42752: data = 8'hf9;
      17'd42753: data = 8'h00;
      17'd42754: data = 8'hf9;
      17'd42755: data = 8'hf5;
      17'd42756: data = 8'hf2;
      17'd42757: data = 8'hf6;
      17'd42758: data = 8'hf4;
      17'd42759: data = 8'hf4;
      17'd42760: data = 8'h00;
      17'd42761: data = 8'hf9;
      17'd42762: data = 8'hf1;
      17'd42763: data = 8'hf4;
      17'd42764: data = 8'hfc;
      17'd42765: data = 8'hf9;
      17'd42766: data = 8'hf6;
      17'd42767: data = 8'h00;
      17'd42768: data = 8'hfe;
      17'd42769: data = 8'hf6;
      17'd42770: data = 8'hfe;
      17'd42771: data = 8'hfd;
      17'd42772: data = 8'hed;
      17'd42773: data = 8'hf9;
      17'd42774: data = 8'hfc;
      17'd42775: data = 8'hed;
      17'd42776: data = 8'hf9;
      17'd42777: data = 8'hfc;
      17'd42778: data = 8'hed;
      17'd42779: data = 8'hf6;
      17'd42780: data = 8'hfe;
      17'd42781: data = 8'hf9;
      17'd42782: data = 8'hf1;
      17'd42783: data = 8'hf5;
      17'd42784: data = 8'hf6;
      17'd42785: data = 8'hef;
      17'd42786: data = 8'hf4;
      17'd42787: data = 8'hfd;
      17'd42788: data = 8'hf4;
      17'd42789: data = 8'hf1;
      17'd42790: data = 8'hf5;
      17'd42791: data = 8'hf6;
      17'd42792: data = 8'hfa;
      17'd42793: data = 8'hfc;
      17'd42794: data = 8'hf5;
      17'd42795: data = 8'hfe;
      17'd42796: data = 8'hfe;
      17'd42797: data = 8'hf6;
      17'd42798: data = 8'hfa;
      17'd42799: data = 8'hfe;
      17'd42800: data = 8'hf5;
      17'd42801: data = 8'hec;
      17'd42802: data = 8'hfa;
      17'd42803: data = 8'hfa;
      17'd42804: data = 8'hef;
      17'd42805: data = 8'hf6;
      17'd42806: data = 8'hf5;
      17'd42807: data = 8'hf5;
      17'd42808: data = 8'hfe;
      17'd42809: data = 8'hfd;
      17'd42810: data = 8'hf9;
      17'd42811: data = 8'hfe;
      17'd42812: data = 8'hfa;
      17'd42813: data = 8'hf9;
      17'd42814: data = 8'h00;
      17'd42815: data = 8'hfe;
      17'd42816: data = 8'hef;
      17'd42817: data = 8'hf2;
      17'd42818: data = 8'hfa;
      17'd42819: data = 8'hf9;
      17'd42820: data = 8'hf5;
      17'd42821: data = 8'hf9;
      17'd42822: data = 8'hf9;
      17'd42823: data = 8'hf4;
      17'd42824: data = 8'hfe;
      17'd42825: data = 8'h02;
      17'd42826: data = 8'hfd;
      17'd42827: data = 8'hfa;
      17'd42828: data = 8'hfd;
      17'd42829: data = 8'hfe;
      17'd42830: data = 8'hfd;
      17'd42831: data = 8'hfd;
      17'd42832: data = 8'hfa;
      17'd42833: data = 8'hf9;
      17'd42834: data = 8'hfe;
      17'd42835: data = 8'hfc;
      17'd42836: data = 8'hfa;
      17'd42837: data = 8'h00;
      17'd42838: data = 8'hfa;
      17'd42839: data = 8'hfa;
      17'd42840: data = 8'h00;
      17'd42841: data = 8'hfa;
      17'd42842: data = 8'hfc;
      17'd42843: data = 8'hfc;
      17'd42844: data = 8'hfd;
      17'd42845: data = 8'hfa;
      17'd42846: data = 8'hf6;
      17'd42847: data = 8'hfa;
      17'd42848: data = 8'hfc;
      17'd42849: data = 8'hfc;
      17'd42850: data = 8'hfc;
      17'd42851: data = 8'hfc;
      17'd42852: data = 8'hfd;
      17'd42853: data = 8'h04;
      17'd42854: data = 8'h06;
      17'd42855: data = 8'h01;
      17'd42856: data = 8'h01;
      17'd42857: data = 8'h02;
      17'd42858: data = 8'h00;
      17'd42859: data = 8'hfe;
      17'd42860: data = 8'h02;
      17'd42861: data = 8'hfe;
      17'd42862: data = 8'hfe;
      17'd42863: data = 8'h02;
      17'd42864: data = 8'h05;
      17'd42865: data = 8'h05;
      17'd42866: data = 8'h02;
      17'd42867: data = 8'h01;
      17'd42868: data = 8'h09;
      17'd42869: data = 8'h0a;
      17'd42870: data = 8'h06;
      17'd42871: data = 8'h06;
      17'd42872: data = 8'h05;
      17'd42873: data = 8'h02;
      17'd42874: data = 8'h01;
      17'd42875: data = 8'h05;
      17'd42876: data = 8'h01;
      17'd42877: data = 8'h00;
      17'd42878: data = 8'h04;
      17'd42879: data = 8'h00;
      17'd42880: data = 8'h01;
      17'd42881: data = 8'h0a;
      17'd42882: data = 8'h06;
      17'd42883: data = 8'h04;
      17'd42884: data = 8'h0a;
      17'd42885: data = 8'h09;
      17'd42886: data = 8'h05;
      17'd42887: data = 8'h06;
      17'd42888: data = 8'h0d;
      17'd42889: data = 8'h04;
      17'd42890: data = 8'h00;
      17'd42891: data = 8'h06;
      17'd42892: data = 8'h00;
      17'd42893: data = 8'hfd;
      17'd42894: data = 8'h00;
      17'd42895: data = 8'h01;
      17'd42896: data = 8'h00;
      17'd42897: data = 8'h04;
      17'd42898: data = 8'h0c;
      17'd42899: data = 8'h06;
      17'd42900: data = 8'h06;
      17'd42901: data = 8'h0c;
      17'd42902: data = 8'h0a;
      17'd42903: data = 8'h0a;
      17'd42904: data = 8'h0c;
      17'd42905: data = 8'h06;
      17'd42906: data = 8'h06;
      17'd42907: data = 8'h09;
      17'd42908: data = 8'h05;
      17'd42909: data = 8'h04;
      17'd42910: data = 8'h04;
      17'd42911: data = 8'h06;
      17'd42912: data = 8'h01;
      17'd42913: data = 8'h02;
      17'd42914: data = 8'h06;
      17'd42915: data = 8'h04;
      17'd42916: data = 8'h09;
      17'd42917: data = 8'h0c;
      17'd42918: data = 8'h09;
      17'd42919: data = 8'h06;
      17'd42920: data = 8'h06;
      17'd42921: data = 8'h05;
      17'd42922: data = 8'h01;
      17'd42923: data = 8'h04;
      17'd42924: data = 8'h04;
      17'd42925: data = 8'h00;
      17'd42926: data = 8'h02;
      17'd42927: data = 8'h02;
      17'd42928: data = 8'h01;
      17'd42929: data = 8'h05;
      17'd42930: data = 8'h06;
      17'd42931: data = 8'h04;
      17'd42932: data = 8'h04;
      17'd42933: data = 8'h06;
      17'd42934: data = 8'h05;
      17'd42935: data = 8'h06;
      17'd42936: data = 8'h09;
      17'd42937: data = 8'h05;
      17'd42938: data = 8'h04;
      17'd42939: data = 8'h01;
      17'd42940: data = 8'h00;
      17'd42941: data = 8'h02;
      17'd42942: data = 8'h02;
      17'd42943: data = 8'h00;
      17'd42944: data = 8'hfe;
      17'd42945: data = 8'h04;
      17'd42946: data = 8'h05;
      17'd42947: data = 8'h04;
      17'd42948: data = 8'h04;
      17'd42949: data = 8'h06;
      17'd42950: data = 8'h06;
      17'd42951: data = 8'h05;
      17'd42952: data = 8'h05;
      17'd42953: data = 8'h05;
      17'd42954: data = 8'h05;
      17'd42955: data = 8'h06;
      17'd42956: data = 8'h05;
      17'd42957: data = 8'h04;
      17'd42958: data = 8'h04;
      17'd42959: data = 8'h04;
      17'd42960: data = 8'h02;
      17'd42961: data = 8'h02;
      17'd42962: data = 8'h05;
      17'd42963: data = 8'h04;
      17'd42964: data = 8'h04;
      17'd42965: data = 8'h05;
      17'd42966: data = 8'h02;
      17'd42967: data = 8'h01;
      17'd42968: data = 8'h02;
      17'd42969: data = 8'h04;
      17'd42970: data = 8'h01;
      17'd42971: data = 8'h00;
      17'd42972: data = 8'h00;
      17'd42973: data = 8'h00;
      17'd42974: data = 8'h05;
      17'd42975: data = 8'h05;
      17'd42976: data = 8'h00;
      17'd42977: data = 8'h00;
      17'd42978: data = 8'h00;
      17'd42979: data = 8'h01;
      17'd42980: data = 8'h02;
      17'd42981: data = 8'h00;
      17'd42982: data = 8'hfe;
      17'd42983: data = 8'h01;
      17'd42984: data = 8'h02;
      17'd42985: data = 8'h02;
      17'd42986: data = 8'h00;
      17'd42987: data = 8'hfe;
      17'd42988: data = 8'hfe;
      17'd42989: data = 8'hfe;
      17'd42990: data = 8'h00;
      17'd42991: data = 8'h02;
      17'd42992: data = 8'h00;
      17'd42993: data = 8'hfe;
      17'd42994: data = 8'h00;
      17'd42995: data = 8'h01;
      17'd42996: data = 8'h00;
      17'd42997: data = 8'h00;
      17'd42998: data = 8'h00;
      17'd42999: data = 8'hfd;
      17'd43000: data = 8'hfe;
      17'd43001: data = 8'h00;
      17'd43002: data = 8'h01;
      17'd43003: data = 8'hfe;
      17'd43004: data = 8'hfc;
      17'd43005: data = 8'hfe;
      17'd43006: data = 8'h01;
      17'd43007: data = 8'h02;
      17'd43008: data = 8'h01;
      17'd43009: data = 8'hfc;
      17'd43010: data = 8'hfe;
      17'd43011: data = 8'h01;
      17'd43012: data = 8'hfe;
      17'd43013: data = 8'hfd;
      17'd43014: data = 8'hfe;
      17'd43015: data = 8'hfe;
      17'd43016: data = 8'hfc;
      17'd43017: data = 8'hfe;
      17'd43018: data = 8'h00;
      17'd43019: data = 8'hfd;
      17'd43020: data = 8'hfd;
      17'd43021: data = 8'h00;
      17'd43022: data = 8'h01;
      17'd43023: data = 8'hfd;
      17'd43024: data = 8'hfa;
      17'd43025: data = 8'hfa;
      17'd43026: data = 8'hfd;
      17'd43027: data = 8'hfd;
      17'd43028: data = 8'hfc;
      17'd43029: data = 8'hfa;
      17'd43030: data = 8'hfc;
      17'd43031: data = 8'h00;
      17'd43032: data = 8'h00;
      17'd43033: data = 8'h00;
      17'd43034: data = 8'hfe;
      17'd43035: data = 8'h00;
      17'd43036: data = 8'h00;
      17'd43037: data = 8'hfd;
      17'd43038: data = 8'hfc;
      17'd43039: data = 8'hfd;
      17'd43040: data = 8'h00;
      17'd43041: data = 8'hfd;
      17'd43042: data = 8'hfd;
      17'd43043: data = 8'hfd;
      17'd43044: data = 8'hfc;
      17'd43045: data = 8'hfd;
      17'd43046: data = 8'h01;
      17'd43047: data = 8'h01;
      17'd43048: data = 8'h00;
      17'd43049: data = 8'h02;
      17'd43050: data = 8'h01;
      17'd43051: data = 8'hfd;
      17'd43052: data = 8'h00;
      17'd43053: data = 8'h00;
      17'd43054: data = 8'hfa;
      17'd43055: data = 8'hfd;
      17'd43056: data = 8'hfd;
      17'd43057: data = 8'hfa;
      17'd43058: data = 8'hfd;
      17'd43059: data = 8'h00;
      17'd43060: data = 8'hfd;
      17'd43061: data = 8'hf9;
      17'd43062: data = 8'h01;
      17'd43063: data = 8'hfe;
      17'd43064: data = 8'hf9;
      17'd43065: data = 8'hfe;
      17'd43066: data = 8'hfe;
      17'd43067: data = 8'hf9;
      17'd43068: data = 8'hfc;
      17'd43069: data = 8'hfd;
      17'd43070: data = 8'hfc;
      17'd43071: data = 8'hf9;
      17'd43072: data = 8'hfa;
      17'd43073: data = 8'hfd;
      17'd43074: data = 8'hfc;
      17'd43075: data = 8'hfa;
      17'd43076: data = 8'hfc;
      17'd43077: data = 8'hf9;
      17'd43078: data = 8'hf5;
      17'd43079: data = 8'hfc;
      17'd43080: data = 8'hfc;
      17'd43081: data = 8'hf2;
      17'd43082: data = 8'hf6;
      17'd43083: data = 8'hfa;
      17'd43084: data = 8'hf6;
      17'd43085: data = 8'hfd;
      17'd43086: data = 8'hfd;
      17'd43087: data = 8'hfc;
      17'd43088: data = 8'hfc;
      17'd43089: data = 8'hf9;
      17'd43090: data = 8'hf9;
      17'd43091: data = 8'hf9;
      17'd43092: data = 8'hf6;
      17'd43093: data = 8'hfa;
      17'd43094: data = 8'hfc;
      17'd43095: data = 8'hfa;
      17'd43096: data = 8'hfc;
      17'd43097: data = 8'hf9;
      17'd43098: data = 8'hfd;
      17'd43099: data = 8'hfc;
      17'd43100: data = 8'hfa;
      17'd43101: data = 8'h00;
      17'd43102: data = 8'hfe;
      17'd43103: data = 8'hfc;
      17'd43104: data = 8'hfd;
      17'd43105: data = 8'h01;
      17'd43106: data = 8'h00;
      17'd43107: data = 8'hfc;
      17'd43108: data = 8'hfe;
      17'd43109: data = 8'hfa;
      17'd43110: data = 8'hf6;
      17'd43111: data = 8'hf9;
      17'd43112: data = 8'hfa;
      17'd43113: data = 8'hfc;
      17'd43114: data = 8'hfc;
      17'd43115: data = 8'h01;
      17'd43116: data = 8'hfe;
      17'd43117: data = 8'hf6;
      17'd43118: data = 8'hfe;
      17'd43119: data = 8'hfd;
      17'd43120: data = 8'hf6;
      17'd43121: data = 8'hfe;
      17'd43122: data = 8'hfd;
      17'd43123: data = 8'hfa;
      17'd43124: data = 8'hfa;
      17'd43125: data = 8'hf9;
      17'd43126: data = 8'hfc;
      17'd43127: data = 8'hfc;
      17'd43128: data = 8'hf9;
      17'd43129: data = 8'hf5;
      17'd43130: data = 8'hf9;
      17'd43131: data = 8'hfc;
      17'd43132: data = 8'hf6;
      17'd43133: data = 8'hf6;
      17'd43134: data = 8'h00;
      17'd43135: data = 8'h00;
      17'd43136: data = 8'hfa;
      17'd43137: data = 8'hf9;
      17'd43138: data = 8'hfd;
      17'd43139: data = 8'hfd;
      17'd43140: data = 8'hfc;
      17'd43141: data = 8'h01;
      17'd43142: data = 8'hfd;
      17'd43143: data = 8'hf6;
      17'd43144: data = 8'hfc;
      17'd43145: data = 8'hfe;
      17'd43146: data = 8'h00;
      17'd43147: data = 8'hfe;
      17'd43148: data = 8'hfc;
      17'd43149: data = 8'hfa;
      17'd43150: data = 8'h00;
      17'd43151: data = 8'h05;
      17'd43152: data = 8'h04;
      17'd43153: data = 8'hfe;
      17'd43154: data = 8'h00;
      17'd43155: data = 8'hfd;
      17'd43156: data = 8'hfd;
      17'd43157: data = 8'h04;
      17'd43158: data = 8'h00;
      17'd43159: data = 8'hf9;
      17'd43160: data = 8'hf9;
      17'd43161: data = 8'h02;
      17'd43162: data = 8'h02;
      17'd43163: data = 8'hfc;
      17'd43164: data = 8'h01;
      17'd43165: data = 8'h00;
      17'd43166: data = 8'h00;
      17'd43167: data = 8'h05;
      17'd43168: data = 8'h04;
      17'd43169: data = 8'h01;
      17'd43170: data = 8'h02;
      17'd43171: data = 8'h05;
      17'd43172: data = 8'h01;
      17'd43173: data = 8'h02;
      17'd43174: data = 8'h04;
      17'd43175: data = 8'hfe;
      17'd43176: data = 8'hfc;
      17'd43177: data = 8'h00;
      17'd43178: data = 8'h05;
      17'd43179: data = 8'h00;
      17'd43180: data = 8'h00;
      17'd43181: data = 8'h05;
      17'd43182: data = 8'h01;
      17'd43183: data = 8'hfe;
      17'd43184: data = 8'h04;
      17'd43185: data = 8'h02;
      17'd43186: data = 8'h00;
      17'd43187: data = 8'h01;
      17'd43188: data = 8'h02;
      17'd43189: data = 8'h04;
      17'd43190: data = 8'h05;
      17'd43191: data = 8'h06;
      17'd43192: data = 8'h02;
      17'd43193: data = 8'h04;
      17'd43194: data = 8'h01;
      17'd43195: data = 8'h02;
      17'd43196: data = 8'h04;
      17'd43197: data = 8'h05;
      17'd43198: data = 8'h01;
      17'd43199: data = 8'h01;
      17'd43200: data = 8'h06;
      17'd43201: data = 8'h02;
      17'd43202: data = 8'h02;
      17'd43203: data = 8'h09;
      17'd43204: data = 8'h04;
      17'd43205: data = 8'h00;
      17'd43206: data = 8'h04;
      17'd43207: data = 8'h0a;
      17'd43208: data = 8'h05;
      17'd43209: data = 8'h06;
      17'd43210: data = 8'h05;
      17'd43211: data = 8'h01;
      17'd43212: data = 8'hfe;
      17'd43213: data = 8'h01;
      17'd43214: data = 8'h01;
      17'd43215: data = 8'h00;
      17'd43216: data = 8'h02;
      17'd43217: data = 8'h01;
      17'd43218: data = 8'h04;
      17'd43219: data = 8'h09;
      17'd43220: data = 8'h09;
      17'd43221: data = 8'h05;
      17'd43222: data = 8'h06;
      17'd43223: data = 8'h06;
      17'd43224: data = 8'h05;
      17'd43225: data = 8'h05;
      17'd43226: data = 8'h05;
      17'd43227: data = 8'h04;
      17'd43228: data = 8'h01;
      17'd43229: data = 8'h01;
      17'd43230: data = 8'h02;
      17'd43231: data = 8'h01;
      17'd43232: data = 8'hfe;
      17'd43233: data = 8'h05;
      17'd43234: data = 8'h02;
      17'd43235: data = 8'h01;
      17'd43236: data = 8'h06;
      17'd43237: data = 8'h04;
      17'd43238: data = 8'h04;
      17'd43239: data = 8'h02;
      17'd43240: data = 8'hfe;
      17'd43241: data = 8'hfe;
      17'd43242: data = 8'h02;
      17'd43243: data = 8'h01;
      17'd43244: data = 8'hfd;
      17'd43245: data = 8'h01;
      17'd43246: data = 8'h01;
      17'd43247: data = 8'hfe;
      17'd43248: data = 8'h01;
      17'd43249: data = 8'h05;
      17'd43250: data = 8'h04;
      17'd43251: data = 8'h02;
      17'd43252: data = 8'h05;
      17'd43253: data = 8'h0a;
      17'd43254: data = 8'h09;
      17'd43255: data = 8'h04;
      17'd43256: data = 8'h06;
      17'd43257: data = 8'h05;
      17'd43258: data = 8'h02;
      17'd43259: data = 8'h02;
      17'd43260: data = 8'h04;
      17'd43261: data = 8'h01;
      17'd43262: data = 8'hfe;
      17'd43263: data = 8'hfe;
      17'd43264: data = 8'hfe;
      17'd43265: data = 8'hfe;
      17'd43266: data = 8'hfe;
      17'd43267: data = 8'h00;
      17'd43268: data = 8'hfe;
      17'd43269: data = 8'h00;
      17'd43270: data = 8'h00;
      17'd43271: data = 8'h01;
      17'd43272: data = 8'h02;
      17'd43273: data = 8'h00;
      17'd43274: data = 8'h00;
      17'd43275: data = 8'h01;
      17'd43276: data = 8'h01;
      17'd43277: data = 8'hfe;
      17'd43278: data = 8'hfd;
      17'd43279: data = 8'h00;
      17'd43280: data = 8'hfe;
      17'd43281: data = 8'hfe;
      17'd43282: data = 8'h02;
      17'd43283: data = 8'h01;
      17'd43284: data = 8'hfe;
      17'd43285: data = 8'hfd;
      17'd43286: data = 8'h01;
      17'd43287: data = 8'h00;
      17'd43288: data = 8'hfe;
      17'd43289: data = 8'hfd;
      17'd43290: data = 8'hfc;
      17'd43291: data = 8'h01;
      17'd43292: data = 8'hfe;
      17'd43293: data = 8'hfd;
      17'd43294: data = 8'hfe;
      17'd43295: data = 8'hfc;
      17'd43296: data = 8'hfa;
      17'd43297: data = 8'h00;
      17'd43298: data = 8'h02;
      17'd43299: data = 8'h01;
      17'd43300: data = 8'h00;
      17'd43301: data = 8'h01;
      17'd43302: data = 8'h02;
      17'd43303: data = 8'h04;
      17'd43304: data = 8'hfd;
      17'd43305: data = 8'hfe;
      17'd43306: data = 8'h01;
      17'd43307: data = 8'h00;
      17'd43308: data = 8'h00;
      17'd43309: data = 8'h01;
      17'd43310: data = 8'h02;
      17'd43311: data = 8'h01;
      17'd43312: data = 8'h01;
      17'd43313: data = 8'hfd;
      17'd43314: data = 8'hfe;
      17'd43315: data = 8'h00;
      17'd43316: data = 8'hfd;
      17'd43317: data = 8'hfd;
      17'd43318: data = 8'hfe;
      17'd43319: data = 8'hfe;
      17'd43320: data = 8'hfc;
      17'd43321: data = 8'hfc;
      17'd43322: data = 8'hfc;
      17'd43323: data = 8'hfa;
      17'd43324: data = 8'hfc;
      17'd43325: data = 8'hfc;
      17'd43326: data = 8'hfc;
      17'd43327: data = 8'hfd;
      17'd43328: data = 8'hfd;
      17'd43329: data = 8'hfd;
      17'd43330: data = 8'hfe;
      17'd43331: data = 8'hfc;
      17'd43332: data = 8'hfc;
      17'd43333: data = 8'hfd;
      17'd43334: data = 8'hfd;
      17'd43335: data = 8'hfa;
      17'd43336: data = 8'hf9;
      17'd43337: data = 8'hfa;
      17'd43338: data = 8'hfa;
      17'd43339: data = 8'hf9;
      17'd43340: data = 8'hfa;
      17'd43341: data = 8'hfa;
      17'd43342: data = 8'hfc;
      17'd43343: data = 8'hfd;
      17'd43344: data = 8'hfd;
      17'd43345: data = 8'hfd;
      17'd43346: data = 8'hfd;
      17'd43347: data = 8'hfc;
      17'd43348: data = 8'h00;
      17'd43349: data = 8'h01;
      17'd43350: data = 8'hfd;
      17'd43351: data = 8'hfd;
      17'd43352: data = 8'hfc;
      17'd43353: data = 8'hfd;
      17'd43354: data = 8'h00;
      17'd43355: data = 8'hfd;
      17'd43356: data = 8'hfc;
      17'd43357: data = 8'hfe;
      17'd43358: data = 8'hfe;
      17'd43359: data = 8'hfe;
      17'd43360: data = 8'hfe;
      17'd43361: data = 8'hfe;
      17'd43362: data = 8'hfe;
      17'd43363: data = 8'hfd;
      17'd43364: data = 8'hfd;
      17'd43365: data = 8'hfe;
      17'd43366: data = 8'hfc;
      17'd43367: data = 8'hfc;
      17'd43368: data = 8'hfc;
      17'd43369: data = 8'hfc;
      17'd43370: data = 8'hfc;
      17'd43371: data = 8'hfa;
      17'd43372: data = 8'hfc;
      17'd43373: data = 8'hfa;
      17'd43374: data = 8'hfc;
      17'd43375: data = 8'hfc;
      17'd43376: data = 8'hfa;
      17'd43377: data = 8'hfa;
      17'd43378: data = 8'hfe;
      17'd43379: data = 8'hfe;
      17'd43380: data = 8'hfa;
      17'd43381: data = 8'hfa;
      17'd43382: data = 8'hfc;
      17'd43383: data = 8'hfc;
      17'd43384: data = 8'hfc;
      17'd43385: data = 8'hfc;
      17'd43386: data = 8'hf9;
      17'd43387: data = 8'hfa;
      17'd43388: data = 8'hfa;
      17'd43389: data = 8'hfa;
      17'd43390: data = 8'hfa;
      17'd43391: data = 8'hfa;
      17'd43392: data = 8'hf9;
      17'd43393: data = 8'hf9;
      17'd43394: data = 8'hfc;
      17'd43395: data = 8'hfe;
      17'd43396: data = 8'hfa;
      17'd43397: data = 8'hfa;
      17'd43398: data = 8'hfa;
      17'd43399: data = 8'hfc;
      17'd43400: data = 8'hfc;
      17'd43401: data = 8'hfa;
      17'd43402: data = 8'hfa;
      17'd43403: data = 8'hfc;
      17'd43404: data = 8'hfc;
      17'd43405: data = 8'hfa;
      17'd43406: data = 8'hfe;
      17'd43407: data = 8'hfe;
      17'd43408: data = 8'hfd;
      17'd43409: data = 8'hfc;
      17'd43410: data = 8'hfd;
      17'd43411: data = 8'hfd;
      17'd43412: data = 8'hfe;
      17'd43413: data = 8'hfd;
      17'd43414: data = 8'hfc;
      17'd43415: data = 8'hfe;
      17'd43416: data = 8'hfe;
      17'd43417: data = 8'hfe;
      17'd43418: data = 8'hfd;
      17'd43419: data = 8'hfe;
      17'd43420: data = 8'hfe;
      17'd43421: data = 8'hfd;
      17'd43422: data = 8'hfd;
      17'd43423: data = 8'hfe;
      17'd43424: data = 8'hfd;
      17'd43425: data = 8'hfd;
      17'd43426: data = 8'hfc;
      17'd43427: data = 8'hfc;
      17'd43428: data = 8'hfa;
      17'd43429: data = 8'hf9;
      17'd43430: data = 8'hfc;
      17'd43431: data = 8'hfd;
      17'd43432: data = 8'hfd;
      17'd43433: data = 8'hfd;
      17'd43434: data = 8'hfc;
      17'd43435: data = 8'hfe;
      17'd43436: data = 8'h01;
      17'd43437: data = 8'h01;
      17'd43438: data = 8'h01;
      17'd43439: data = 8'h00;
      17'd43440: data = 8'h00;
      17'd43441: data = 8'h01;
      17'd43442: data = 8'h00;
      17'd43443: data = 8'h00;
      17'd43444: data = 8'hfe;
      17'd43445: data = 8'h00;
      17'd43446: data = 8'h01;
      17'd43447: data = 8'hfe;
      17'd43448: data = 8'hfe;
      17'd43449: data = 8'h00;
      17'd43450: data = 8'h01;
      17'd43451: data = 8'h00;
      17'd43452: data = 8'h00;
      17'd43453: data = 8'h00;
      17'd43454: data = 8'h01;
      17'd43455: data = 8'h04;
      17'd43456: data = 8'h05;
      17'd43457: data = 8'h02;
      17'd43458: data = 8'h00;
      17'd43459: data = 8'h02;
      17'd43460: data = 8'h04;
      17'd43461: data = 8'h05;
      17'd43462: data = 8'h01;
      17'd43463: data = 8'h01;
      17'd43464: data = 8'h01;
      17'd43465: data = 8'h02;
      17'd43466: data = 8'h05;
      17'd43467: data = 8'h02;
      17'd43468: data = 8'h05;
      17'd43469: data = 8'h05;
      17'd43470: data = 8'h05;
      17'd43471: data = 8'h06;
      17'd43472: data = 8'h04;
      17'd43473: data = 8'h04;
      17'd43474: data = 8'h04;
      17'd43475: data = 8'h04;
      17'd43476: data = 8'h02;
      17'd43477: data = 8'h01;
      17'd43478: data = 8'h00;
      17'd43479: data = 8'hfe;
      17'd43480: data = 8'h00;
      17'd43481: data = 8'h02;
      17'd43482: data = 8'h02;
      17'd43483: data = 8'h01;
      17'd43484: data = 8'h02;
      17'd43485: data = 8'h05;
      17'd43486: data = 8'h02;
      17'd43487: data = 8'h01;
      17'd43488: data = 8'h04;
      17'd43489: data = 8'h04;
      17'd43490: data = 8'h01;
      17'd43491: data = 8'h02;
      17'd43492: data = 8'h04;
      17'd43493: data = 8'h01;
      17'd43494: data = 8'h04;
      17'd43495: data = 8'h04;
      17'd43496: data = 8'h01;
      17'd43497: data = 8'h01;
      17'd43498: data = 8'h01;
      17'd43499: data = 8'h04;
      17'd43500: data = 8'h01;
      17'd43501: data = 8'h02;
      17'd43502: data = 8'h02;
      17'd43503: data = 8'h00;
      17'd43504: data = 8'hfe;
      17'd43505: data = 8'hfe;
      17'd43506: data = 8'hfd;
      17'd43507: data = 8'hfd;
      17'd43508: data = 8'h00;
      17'd43509: data = 8'h00;
      17'd43510: data = 8'h01;
      17'd43511: data = 8'h01;
      17'd43512: data = 8'h01;
      17'd43513: data = 8'h02;
      17'd43514: data = 8'h00;
      17'd43515: data = 8'h01;
      17'd43516: data = 8'h00;
      17'd43517: data = 8'hfd;
      17'd43518: data = 8'h01;
      17'd43519: data = 8'h01;
      17'd43520: data = 8'h00;
      17'd43521: data = 8'h00;
      17'd43522: data = 8'h01;
      17'd43523: data = 8'h01;
      17'd43524: data = 8'h01;
      17'd43525: data = 8'h02;
      17'd43526: data = 8'h01;
      17'd43527: data = 8'h00;
      17'd43528: data = 8'h01;
      17'd43529: data = 8'h02;
      17'd43530: data = 8'hfe;
      17'd43531: data = 8'hfd;
      17'd43532: data = 8'h00;
      17'd43533: data = 8'h00;
      17'd43534: data = 8'hfe;
      17'd43535: data = 8'hfe;
      17'd43536: data = 8'hfe;
      17'd43537: data = 8'hfe;
      17'd43538: data = 8'h01;
      17'd43539: data = 8'h01;
      17'd43540: data = 8'h01;
      17'd43541: data = 8'hfe;
      17'd43542: data = 8'h00;
      17'd43543: data = 8'h02;
      17'd43544: data = 8'h01;
      17'd43545: data = 8'h02;
      17'd43546: data = 8'h01;
      17'd43547: data = 8'hfe;
      17'd43548: data = 8'h00;
      17'd43549: data = 8'h00;
      17'd43550: data = 8'hfe;
      17'd43551: data = 8'hfe;
      17'd43552: data = 8'h00;
      17'd43553: data = 8'h00;
      17'd43554: data = 8'h00;
      17'd43555: data = 8'h00;
      17'd43556: data = 8'h00;
      17'd43557: data = 8'h00;
      17'd43558: data = 8'h00;
      17'd43559: data = 8'hfe;
      17'd43560: data = 8'hfd;
      17'd43561: data = 8'hfe;
      17'd43562: data = 8'hfe;
      17'd43563: data = 8'h00;
      17'd43564: data = 8'hfe;
      17'd43565: data = 8'hfe;
      17'd43566: data = 8'h00;
      17'd43567: data = 8'h00;
      17'd43568: data = 8'h01;
      17'd43569: data = 8'h00;
      17'd43570: data = 8'hfd;
      17'd43571: data = 8'hfd;
      17'd43572: data = 8'hfd;
      17'd43573: data = 8'hfd;
      17'd43574: data = 8'hfe;
      17'd43575: data = 8'hfd;
      17'd43576: data = 8'hfd;
      17'd43577: data = 8'hfd;
      17'd43578: data = 8'hfd;
      17'd43579: data = 8'h00;
      17'd43580: data = 8'hfd;
      17'd43581: data = 8'hfe;
      17'd43582: data = 8'hfe;
      17'd43583: data = 8'h00;
      17'd43584: data = 8'h01;
      17'd43585: data = 8'h00;
      17'd43586: data = 8'h00;
      17'd43587: data = 8'h00;
      17'd43588: data = 8'h01;
      17'd43589: data = 8'h01;
      17'd43590: data = 8'hfe;
      17'd43591: data = 8'hfd;
      17'd43592: data = 8'h00;
      17'd43593: data = 8'h00;
      17'd43594: data = 8'hfd;
      17'd43595: data = 8'h00;
      17'd43596: data = 8'h00;
      17'd43597: data = 8'hfe;
      17'd43598: data = 8'h00;
      17'd43599: data = 8'hfe;
      17'd43600: data = 8'hfd;
      17'd43601: data = 8'hfe;
      17'd43602: data = 8'hfc;
      17'd43603: data = 8'hfc;
      17'd43604: data = 8'hfe;
      17'd43605: data = 8'hfe;
      17'd43606: data = 8'hfc;
      17'd43607: data = 8'hfa;
      17'd43608: data = 8'hfc;
      17'd43609: data = 8'hfc;
      17'd43610: data = 8'hfa;
      17'd43611: data = 8'hfa;
      17'd43612: data = 8'hfd;
      17'd43613: data = 8'hfd;
      17'd43614: data = 8'hfc;
      17'd43615: data = 8'h00;
      17'd43616: data = 8'h00;
      17'd43617: data = 8'hfe;
      17'd43618: data = 8'h01;
      17'd43619: data = 8'h00;
      17'd43620: data = 8'hfe;
      17'd43621: data = 8'h00;
      17'd43622: data = 8'h00;
      17'd43623: data = 8'hfe;
      17'd43624: data = 8'hfd;
      17'd43625: data = 8'hfd;
      17'd43626: data = 8'hfd;
      17'd43627: data = 8'hfd;
      17'd43628: data = 8'hfa;
      17'd43629: data = 8'hfc;
      17'd43630: data = 8'hfd;
      17'd43631: data = 8'hfc;
      17'd43632: data = 8'hfe;
      17'd43633: data = 8'h00;
      17'd43634: data = 8'h00;
      17'd43635: data = 8'h01;
      17'd43636: data = 8'h02;
      17'd43637: data = 8'hfe;
      17'd43638: data = 8'hfe;
      17'd43639: data = 8'hfe;
      17'd43640: data = 8'hfd;
      17'd43641: data = 8'hfe;
      17'd43642: data = 8'hfd;
      17'd43643: data = 8'hfc;
      17'd43644: data = 8'hfc;
      17'd43645: data = 8'hfd;
      17'd43646: data = 8'hfe;
      17'd43647: data = 8'hfd;
      17'd43648: data = 8'hfe;
      17'd43649: data = 8'h01;
      17'd43650: data = 8'h01;
      17'd43651: data = 8'h02;
      17'd43652: data = 8'h01;
      17'd43653: data = 8'h01;
      17'd43654: data = 8'h01;
      17'd43655: data = 8'h01;
      17'd43656: data = 8'h01;
      17'd43657: data = 8'h00;
      17'd43658: data = 8'hfd;
      17'd43659: data = 8'hfe;
      17'd43660: data = 8'h01;
      17'd43661: data = 8'hfe;
      17'd43662: data = 8'hfd;
      17'd43663: data = 8'hfd;
      17'd43664: data = 8'hfe;
      17'd43665: data = 8'h00;
      17'd43666: data = 8'hfe;
      17'd43667: data = 8'hfd;
      17'd43668: data = 8'hfe;
      17'd43669: data = 8'hfe;
      17'd43670: data = 8'h00;
      17'd43671: data = 8'hfe;
      17'd43672: data = 8'hfe;
      17'd43673: data = 8'h00;
      17'd43674: data = 8'hfe;
      17'd43675: data = 8'hfe;
      17'd43676: data = 8'hfe;
      17'd43677: data = 8'hfe;
      17'd43678: data = 8'hfe;
      17'd43679: data = 8'hfc;
      17'd43680: data = 8'hfc;
      17'd43681: data = 8'hfe;
      17'd43682: data = 8'hfe;
      17'd43683: data = 8'hfe;
      17'd43684: data = 8'hfe;
      17'd43685: data = 8'hfd;
      17'd43686: data = 8'hfd;
      17'd43687: data = 8'hfd;
      17'd43688: data = 8'hfe;
      17'd43689: data = 8'hfd;
      17'd43690: data = 8'hfd;
      17'd43691: data = 8'hfe;
      17'd43692: data = 8'hfe;
      17'd43693: data = 8'h00;
      17'd43694: data = 8'hfc;
      17'd43695: data = 8'hfa;
      17'd43696: data = 8'hfe;
      17'd43697: data = 8'hfd;
      17'd43698: data = 8'hfc;
      17'd43699: data = 8'hfd;
      17'd43700: data = 8'hfd;
      17'd43701: data = 8'hfd;
      17'd43702: data = 8'hfd;
      17'd43703: data = 8'hfe;
      17'd43704: data = 8'hfc;
      17'd43705: data = 8'hf9;
      17'd43706: data = 8'hfe;
      17'd43707: data = 8'h00;
      17'd43708: data = 8'hfe;
      17'd43709: data = 8'h00;
      17'd43710: data = 8'h00;
      17'd43711: data = 8'h00;
      17'd43712: data = 8'h00;
      17'd43713: data = 8'hfe;
      17'd43714: data = 8'hfc;
      17'd43715: data = 8'hfd;
      17'd43716: data = 8'hfe;
      17'd43717: data = 8'hfd;
      17'd43718: data = 8'hfc;
      17'd43719: data = 8'hfc;
      17'd43720: data = 8'hfc;
      17'd43721: data = 8'hfd;
      17'd43722: data = 8'hfd;
      17'd43723: data = 8'hfc;
      17'd43724: data = 8'hfe;
      17'd43725: data = 8'hfe;
      17'd43726: data = 8'h00;
      17'd43727: data = 8'hfe;
      17'd43728: data = 8'hfc;
      17'd43729: data = 8'hfd;
      17'd43730: data = 8'hfe;
      17'd43731: data = 8'hfd;
      17'd43732: data = 8'hfc;
      17'd43733: data = 8'hfc;
      17'd43734: data = 8'hfc;
      17'd43735: data = 8'hfc;
      17'd43736: data = 8'hfd;
      17'd43737: data = 8'hfc;
      17'd43738: data = 8'hfd;
      17'd43739: data = 8'h00;
      17'd43740: data = 8'h02;
      17'd43741: data = 8'h01;
      17'd43742: data = 8'hfe;
      17'd43743: data = 8'h00;
      17'd43744: data = 8'h00;
      17'd43745: data = 8'h01;
      17'd43746: data = 8'h02;
      17'd43747: data = 8'h00;
      17'd43748: data = 8'hfd;
      17'd43749: data = 8'hfe;
      17'd43750: data = 8'h02;
      17'd43751: data = 8'h02;
      17'd43752: data = 8'h00;
      17'd43753: data = 8'hfe;
      17'd43754: data = 8'h00;
      17'd43755: data = 8'h01;
      17'd43756: data = 8'h01;
      17'd43757: data = 8'h01;
      17'd43758: data = 8'hfd;
      17'd43759: data = 8'h00;
      17'd43760: data = 8'h01;
      17'd43761: data = 8'hfe;
      17'd43762: data = 8'h00;
      17'd43763: data = 8'hfe;
      17'd43764: data = 8'hfd;
      17'd43765: data = 8'hfe;
      17'd43766: data = 8'hfe;
      17'd43767: data = 8'hfe;
      17'd43768: data = 8'h00;
      17'd43769: data = 8'h00;
      17'd43770: data = 8'h01;
      17'd43771: data = 8'h01;
      17'd43772: data = 8'hfd;
      17'd43773: data = 8'hfe;
      17'd43774: data = 8'h00;
      17'd43775: data = 8'h00;
      17'd43776: data = 8'hfe;
      17'd43777: data = 8'h00;
      17'd43778: data = 8'hfd;
      17'd43779: data = 8'h00;
      17'd43780: data = 8'h02;
      17'd43781: data = 8'h01;
      17'd43782: data = 8'h01;
      17'd43783: data = 8'h01;
      17'd43784: data = 8'h01;
      17'd43785: data = 8'h02;
      17'd43786: data = 8'h02;
      17'd43787: data = 8'h01;
      17'd43788: data = 8'h01;
      17'd43789: data = 8'h02;
      17'd43790: data = 8'h01;
      17'd43791: data = 8'h00;
      17'd43792: data = 8'h00;
      17'd43793: data = 8'h00;
      17'd43794: data = 8'h01;
      17'd43795: data = 8'h00;
      17'd43796: data = 8'h00;
      17'd43797: data = 8'h02;
      17'd43798: data = 8'h02;
      17'd43799: data = 8'h02;
      17'd43800: data = 8'h00;
      17'd43801: data = 8'h00;
      17'd43802: data = 8'h00;
      17'd43803: data = 8'h01;
      17'd43804: data = 8'h05;
      17'd43805: data = 8'h01;
      17'd43806: data = 8'hfe;
      17'd43807: data = 8'h00;
      17'd43808: data = 8'h01;
      17'd43809: data = 8'h01;
      17'd43810: data = 8'hfe;
      17'd43811: data = 8'hfc;
      17'd43812: data = 8'hfc;
      17'd43813: data = 8'hfd;
      17'd43814: data = 8'h00;
      17'd43815: data = 8'h00;
      17'd43816: data = 8'hfe;
      17'd43817: data = 8'hfd;
      17'd43818: data = 8'hfe;
      17'd43819: data = 8'h01;
      17'd43820: data = 8'h01;
      17'd43821: data = 8'hfd;
      17'd43822: data = 8'hfc;
      17'd43823: data = 8'h00;
      17'd43824: data = 8'h01;
      17'd43825: data = 8'h00;
      17'd43826: data = 8'hfd;
      17'd43827: data = 8'hfe;
      17'd43828: data = 8'hfe;
      17'd43829: data = 8'hfe;
      17'd43830: data = 8'h00;
      17'd43831: data = 8'h01;
      17'd43832: data = 8'hfe;
      17'd43833: data = 8'h01;
      17'd43834: data = 8'h00;
      17'd43835: data = 8'h01;
      17'd43836: data = 8'h04;
      17'd43837: data = 8'h01;
      17'd43838: data = 8'h02;
      17'd43839: data = 8'h02;
      17'd43840: data = 8'h00;
      17'd43841: data = 8'h00;
      17'd43842: data = 8'h01;
      17'd43843: data = 8'h00;
      17'd43844: data = 8'hfe;
      17'd43845: data = 8'hfd;
      17'd43846: data = 8'hfe;
      17'd43847: data = 8'h00;
      17'd43848: data = 8'h00;
      17'd43849: data = 8'h00;
      17'd43850: data = 8'h00;
      17'd43851: data = 8'h00;
      17'd43852: data = 8'h00;
      17'd43853: data = 8'h04;
      17'd43854: data = 8'h04;
      17'd43855: data = 8'h02;
      17'd43856: data = 8'h04;
      17'd43857: data = 8'h05;
      17'd43858: data = 8'h04;
      17'd43859: data = 8'h01;
      17'd43860: data = 8'h00;
      17'd43861: data = 8'h01;
      17'd43862: data = 8'h02;
      17'd43863: data = 8'h01;
      17'd43864: data = 8'h00;
      17'd43865: data = 8'hfe;
      17'd43866: data = 8'hfe;
      17'd43867: data = 8'hfe;
      17'd43868: data = 8'h00;
      17'd43869: data = 8'hfe;
      17'd43870: data = 8'hfa;
      17'd43871: data = 8'hfc;
      17'd43872: data = 8'hfe;
      17'd43873: data = 8'hfe;
      17'd43874: data = 8'hfd;
      17'd43875: data = 8'hfc;
      17'd43876: data = 8'hfc;
      17'd43877: data = 8'hfe;
      17'd43878: data = 8'hfe;
      17'd43879: data = 8'hfe;
      17'd43880: data = 8'hfd;
      17'd43881: data = 8'h00;
      17'd43882: data = 8'h00;
      17'd43883: data = 8'hfe;
      17'd43884: data = 8'hfe;
      17'd43885: data = 8'hfd;
      17'd43886: data = 8'hfe;
      17'd43887: data = 8'hfe;
      17'd43888: data = 8'h02;
      17'd43889: data = 8'h00;
      17'd43890: data = 8'hfd;
      17'd43891: data = 8'hfe;
      17'd43892: data = 8'h00;
      17'd43893: data = 8'h01;
      17'd43894: data = 8'h00;
      17'd43895: data = 8'h00;
      17'd43896: data = 8'hfe;
      17'd43897: data = 8'h01;
      17'd43898: data = 8'h01;
      17'd43899: data = 8'hfe;
      17'd43900: data = 8'hfd;
      17'd43901: data = 8'hfe;
      17'd43902: data = 8'h00;
      17'd43903: data = 8'h00;
      17'd43904: data = 8'h00;
      17'd43905: data = 8'hfe;
      17'd43906: data = 8'h00;
      17'd43907: data = 8'h00;
      17'd43908: data = 8'h01;
      17'd43909: data = 8'h02;
      17'd43910: data = 8'h01;
      17'd43911: data = 8'h01;
      17'd43912: data = 8'h00;
      17'd43913: data = 8'h00;
      17'd43914: data = 8'h01;
      17'd43915: data = 8'h01;
      17'd43916: data = 8'h00;
      17'd43917: data = 8'h00;
      17'd43918: data = 8'h00;
      17'd43919: data = 8'h00;
      17'd43920: data = 8'hfe;
      17'd43921: data = 8'hfe;
      17'd43922: data = 8'h00;
      17'd43923: data = 8'hfc;
      17'd43924: data = 8'hfd;
      17'd43925: data = 8'h00;
      17'd43926: data = 8'hfe;
      17'd43927: data = 8'hfe;
      17'd43928: data = 8'hfd;
      17'd43929: data = 8'hfe;
      17'd43930: data = 8'hfe;
      17'd43931: data = 8'hfd;
      17'd43932: data = 8'hfd;
      17'd43933: data = 8'h00;
      17'd43934: data = 8'hfe;
      17'd43935: data = 8'h00;
      17'd43936: data = 8'h01;
      17'd43937: data = 8'h00;
      17'd43938: data = 8'hfe;
      17'd43939: data = 8'h00;
      17'd43940: data = 8'h00;
      17'd43941: data = 8'hfe;
      17'd43942: data = 8'hfd;
      17'd43943: data = 8'hfc;
      17'd43944: data = 8'hfd;
      17'd43945: data = 8'hfd;
      17'd43946: data = 8'hfc;
      17'd43947: data = 8'hfc;
      17'd43948: data = 8'hfd;
      17'd43949: data = 8'hfd;
      17'd43950: data = 8'hfd;
      17'd43951: data = 8'h00;
      17'd43952: data = 8'h02;
      17'd43953: data = 8'h01;
      17'd43954: data = 8'h00;
      17'd43955: data = 8'h02;
      17'd43956: data = 8'h01;
      17'd43957: data = 8'h01;
      17'd43958: data = 8'h00;
      17'd43959: data = 8'hfc;
      17'd43960: data = 8'hfe;
      17'd43961: data = 8'hfd;
      17'd43962: data = 8'hfc;
      17'd43963: data = 8'hfc;
      17'd43964: data = 8'hfc;
      17'd43965: data = 8'hfd;
      17'd43966: data = 8'hfe;
      17'd43967: data = 8'h00;
      17'd43968: data = 8'hfe;
      17'd43969: data = 8'h02;
      17'd43970: data = 8'h02;
      17'd43971: data = 8'h01;
      17'd43972: data = 8'h01;
      17'd43973: data = 8'h01;
      17'd43974: data = 8'hfe;
      17'd43975: data = 8'hfc;
      17'd43976: data = 8'hfe;
      17'd43977: data = 8'hfe;
      17'd43978: data = 8'hfd;
      17'd43979: data = 8'hfd;
      17'd43980: data = 8'h00;
      17'd43981: data = 8'hfe;
      17'd43982: data = 8'hfe;
      17'd43983: data = 8'h02;
      17'd43984: data = 8'h00;
      17'd43985: data = 8'h01;
      17'd43986: data = 8'h04;
      17'd43987: data = 8'h02;
      17'd43988: data = 8'h01;
      17'd43989: data = 8'hfe;
      17'd43990: data = 8'h00;
      17'd43991: data = 8'h00;
      17'd43992: data = 8'hfe;
      17'd43993: data = 8'h00;
      17'd43994: data = 8'hfd;
      17'd43995: data = 8'hfd;
      17'd43996: data = 8'h01;
      17'd43997: data = 8'h02;
      17'd43998: data = 8'h01;
      17'd43999: data = 8'h00;
      17'd44000: data = 8'h00;
      17'd44001: data = 8'h00;
      17'd44002: data = 8'h01;
      17'd44003: data = 8'h00;
      17'd44004: data = 8'hfe;
      17'd44005: data = 8'h00;
      17'd44006: data = 8'hfd;
      17'd44007: data = 8'hfd;
      17'd44008: data = 8'hfe;
      17'd44009: data = 8'h00;
      17'd44010: data = 8'h00;
      17'd44011: data = 8'h01;
      17'd44012: data = 8'h00;
      17'd44013: data = 8'h00;
      17'd44014: data = 8'h04;
      17'd44015: data = 8'h01;
      17'd44016: data = 8'h00;
      17'd44017: data = 8'hfd;
      17'd44018: data = 8'hfe;
      17'd44019: data = 8'h00;
      17'd44020: data = 8'hfe;
      17'd44021: data = 8'hfd;
      17'd44022: data = 8'hfd;
      17'd44023: data = 8'hfe;
      17'd44024: data = 8'hfe;
      17'd44025: data = 8'h02;
      17'd44026: data = 8'h01;
      17'd44027: data = 8'h00;
      17'd44028: data = 8'h01;
      17'd44029: data = 8'h01;
      17'd44030: data = 8'h02;
      17'd44031: data = 8'h00;
      17'd44032: data = 8'hfe;
      17'd44033: data = 8'h00;
      17'd44034: data = 8'hfe;
      17'd44035: data = 8'h01;
      17'd44036: data = 8'hfd;
      17'd44037: data = 8'hfd;
      17'd44038: data = 8'h00;
      17'd44039: data = 8'h00;
      17'd44040: data = 8'h01;
      17'd44041: data = 8'h01;
      17'd44042: data = 8'h01;
      17'd44043: data = 8'h00;
      17'd44044: data = 8'h02;
      17'd44045: data = 8'h00;
      17'd44046: data = 8'hfe;
      17'd44047: data = 8'hfe;
      17'd44048: data = 8'hfd;
      17'd44049: data = 8'h00;
      17'd44050: data = 8'hfe;
      17'd44051: data = 8'hfd;
      17'd44052: data = 8'hfd;
      17'd44053: data = 8'h00;
      17'd44054: data = 8'h01;
      17'd44055: data = 8'h01;
      17'd44056: data = 8'hfe;
      17'd44057: data = 8'h00;
      17'd44058: data = 8'h00;
      17'd44059: data = 8'h01;
      17'd44060: data = 8'h01;
      17'd44061: data = 8'h00;
      17'd44062: data = 8'hfd;
      17'd44063: data = 8'hfc;
      17'd44064: data = 8'hfd;
      17'd44065: data = 8'h00;
      17'd44066: data = 8'hfe;
      17'd44067: data = 8'hfd;
      17'd44068: data = 8'h00;
      17'd44069: data = 8'h00;
      17'd44070: data = 8'h00;
      17'd44071: data = 8'h01;
      17'd44072: data = 8'h01;
      17'd44073: data = 8'hfe;
      17'd44074: data = 8'h01;
      17'd44075: data = 8'h02;
      17'd44076: data = 8'h00;
      17'd44077: data = 8'h02;
      17'd44078: data = 8'h02;
      17'd44079: data = 8'h01;
      17'd44080: data = 8'h02;
      17'd44081: data = 8'h01;
      17'd44082: data = 8'h01;
      17'd44083: data = 8'h01;
      17'd44084: data = 8'h01;
      17'd44085: data = 8'h01;
      17'd44086: data = 8'h00;
      17'd44087: data = 8'h01;
      17'd44088: data = 8'h01;
      17'd44089: data = 8'h01;
      17'd44090: data = 8'hfe;
      17'd44091: data = 8'hfe;
      17'd44092: data = 8'h01;
      17'd44093: data = 8'h02;
      17'd44094: data = 8'h02;
      17'd44095: data = 8'h02;
      17'd44096: data = 8'h02;
      17'd44097: data = 8'h01;
      17'd44098: data = 8'h04;
      17'd44099: data = 8'h04;
      17'd44100: data = 8'h02;
      17'd44101: data = 8'h02;
      17'd44102: data = 8'h02;
      17'd44103: data = 8'h01;
      17'd44104: data = 8'h00;
      17'd44105: data = 8'h00;
      17'd44106: data = 8'hfe;
      17'd44107: data = 8'hfe;
      17'd44108: data = 8'h00;
      17'd44109: data = 8'h01;
      17'd44110: data = 8'hfd;
      17'd44111: data = 8'hfd;
      17'd44112: data = 8'h00;
      17'd44113: data = 8'h01;
      17'd44114: data = 8'h00;
      17'd44115: data = 8'hfd;
      17'd44116: data = 8'hfe;
      17'd44117: data = 8'hfd;
      17'd44118: data = 8'hfe;
      17'd44119: data = 8'hfe;
      17'd44120: data = 8'hfa;
      17'd44121: data = 8'hfd;
      17'd44122: data = 8'hfe;
      17'd44123: data = 8'hfd;
      17'd44124: data = 8'hfd;
      17'd44125: data = 8'hfd;
      17'd44126: data = 8'hfe;
      17'd44127: data = 8'hfd;
      17'd44128: data = 8'h00;
      17'd44129: data = 8'h00;
      17'd44130: data = 8'h00;
      17'd44131: data = 8'h00;
      17'd44132: data = 8'h00;
      17'd44133: data = 8'h01;
      17'd44134: data = 8'hfe;
      17'd44135: data = 8'hfe;
      17'd44136: data = 8'h00;
      17'd44137: data = 8'hfe;
      17'd44138: data = 8'h00;
      17'd44139: data = 8'h00;
      17'd44140: data = 8'h00;
      17'd44141: data = 8'h01;
      17'd44142: data = 8'h00;
      17'd44143: data = 8'h00;
      17'd44144: data = 8'h00;
      17'd44145: data = 8'h00;
      17'd44146: data = 8'h00;
      17'd44147: data = 8'h01;
      17'd44148: data = 8'h02;
      17'd44149: data = 8'h01;
      17'd44150: data = 8'h00;
      17'd44151: data = 8'h01;
      17'd44152: data = 8'h02;
      17'd44153: data = 8'h01;
      17'd44154: data = 8'h02;
      17'd44155: data = 8'h01;
      17'd44156: data = 8'h00;
      17'd44157: data = 8'h01;
      17'd44158: data = 8'h02;
      17'd44159: data = 8'h00;
      17'd44160: data = 8'h00;
      17'd44161: data = 8'hfe;
      17'd44162: data = 8'h00;
      17'd44163: data = 8'hfe;
      17'd44164: data = 8'hfd;
      17'd44165: data = 8'hfd;
      17'd44166: data = 8'hfd;
      17'd44167: data = 8'hfe;
      17'd44168: data = 8'h00;
      17'd44169: data = 8'h00;
      17'd44170: data = 8'hfe;
      17'd44171: data = 8'hfe;
      17'd44172: data = 8'h00;
      17'd44173: data = 8'h01;
      17'd44174: data = 8'h02;
      17'd44175: data = 8'h00;
      17'd44176: data = 8'hfd;
      17'd44177: data = 8'hfe;
      17'd44178: data = 8'h00;
      17'd44179: data = 8'hfe;
      17'd44180: data = 8'hfd;
      17'd44181: data = 8'hfe;
      17'd44182: data = 8'hfe;
      17'd44183: data = 8'hfe;
      17'd44184: data = 8'hfe;
      17'd44185: data = 8'h00;
      17'd44186: data = 8'hfe;
      17'd44187: data = 8'hfe;
      17'd44188: data = 8'h00;
      17'd44189: data = 8'h00;
      17'd44190: data = 8'hfe;
      17'd44191: data = 8'h00;
      17'd44192: data = 8'hfe;
      17'd44193: data = 8'hfd;
      17'd44194: data = 8'hfd;
      17'd44195: data = 8'hfe;
      17'd44196: data = 8'hfe;
      17'd44197: data = 8'hfe;
      17'd44198: data = 8'hfe;
      17'd44199: data = 8'hfd;
      17'd44200: data = 8'hfe;
      17'd44201: data = 8'hfd;
      17'd44202: data = 8'hfd;
      17'd44203: data = 8'hfe;
      17'd44204: data = 8'hfe;
      17'd44205: data = 8'hfd;
      17'd44206: data = 8'hfd;
      17'd44207: data = 8'hfd;
      17'd44208: data = 8'hfe;
      17'd44209: data = 8'h00;
      17'd44210: data = 8'hfe;
      17'd44211: data = 8'hfd;
      17'd44212: data = 8'hfc;
      17'd44213: data = 8'hfd;
      17'd44214: data = 8'h00;
      17'd44215: data = 8'hfc;
      17'd44216: data = 8'hfd;
      17'd44217: data = 8'h01;
      17'd44218: data = 8'h00;
      17'd44219: data = 8'h00;
      17'd44220: data = 8'h00;
      17'd44221: data = 8'h00;
      17'd44222: data = 8'h01;
      17'd44223: data = 8'h00;
      17'd44224: data = 8'hfe;
      17'd44225: data = 8'hfe;
      17'd44226: data = 8'h00;
      17'd44227: data = 8'h00;
      17'd44228: data = 8'hfe;
      17'd44229: data = 8'hfd;
      17'd44230: data = 8'h00;
      17'd44231: data = 8'hfe;
      17'd44232: data = 8'hfe;
      17'd44233: data = 8'h01;
      17'd44234: data = 8'hfe;
      17'd44235: data = 8'hfd;
      17'd44236: data = 8'hfe;
      17'd44237: data = 8'h00;
      17'd44238: data = 8'h00;
      17'd44239: data = 8'h00;
      17'd44240: data = 8'hfe;
      17'd44241: data = 8'hfe;
      17'd44242: data = 8'h00;
      17'd44243: data = 8'h00;
      17'd44244: data = 8'h00;
      17'd44245: data = 8'hfd;
      17'd44246: data = 8'hfd;
      17'd44247: data = 8'hfe;
      17'd44248: data = 8'hfe;
      17'd44249: data = 8'hfe;
      17'd44250: data = 8'hfd;
      17'd44251: data = 8'hfe;
      17'd44252: data = 8'hfe;
      17'd44253: data = 8'h00;
      17'd44254: data = 8'h01;
      17'd44255: data = 8'h00;
      17'd44256: data = 8'hfe;
      17'd44257: data = 8'h00;
      17'd44258: data = 8'h02;
      17'd44259: data = 8'h01;
      17'd44260: data = 8'h00;
      17'd44261: data = 8'hfe;
      17'd44262: data = 8'hfe;
      17'd44263: data = 8'h01;
      17'd44264: data = 8'h00;
      17'd44265: data = 8'hfd;
      17'd44266: data = 8'hfc;
      17'd44267: data = 8'hfd;
      17'd44268: data = 8'h01;
      17'd44269: data = 8'hfe;
      17'd44270: data = 8'hfe;
      17'd44271: data = 8'h00;
      17'd44272: data = 8'h01;
      17'd44273: data = 8'h02;
      17'd44274: data = 8'h01;
      17'd44275: data = 8'h00;
      17'd44276: data = 8'h01;
      17'd44277: data = 8'h01;
      17'd44278: data = 8'h00;
      17'd44279: data = 8'h01;
      17'd44280: data = 8'h02;
      17'd44281: data = 8'h00;
      17'd44282: data = 8'h01;
      17'd44283: data = 8'h00;
      17'd44284: data = 8'hfe;
      17'd44285: data = 8'h00;
      17'd44286: data = 8'h00;
      17'd44287: data = 8'hfc;
      17'd44288: data = 8'hfc;
      17'd44289: data = 8'hfe;
      17'd44290: data = 8'hfe;
      17'd44291: data = 8'h00;
      17'd44292: data = 8'hfe;
      17'd44293: data = 8'hfd;
      17'd44294: data = 8'hfd;
      17'd44295: data = 8'h00;
      17'd44296: data = 8'h01;
      17'd44297: data = 8'h00;
      17'd44298: data = 8'h00;
      17'd44299: data = 8'hfe;
      17'd44300: data = 8'h00;
      17'd44301: data = 8'h01;
      17'd44302: data = 8'h00;
      17'd44303: data = 8'hfd;
      17'd44304: data = 8'hfd;
      17'd44305: data = 8'hfe;
      17'd44306: data = 8'hfe;
      17'd44307: data = 8'hfe;
      17'd44308: data = 8'hfd;
      17'd44309: data = 8'hfd;
      17'd44310: data = 8'hfe;
      17'd44311: data = 8'hfe;
      17'd44312: data = 8'h01;
      17'd44313: data = 8'h00;
      17'd44314: data = 8'hfe;
      17'd44315: data = 8'h00;
      17'd44316: data = 8'h01;
      17'd44317: data = 8'h00;
      17'd44318: data = 8'hfd;
      17'd44319: data = 8'hfe;
      17'd44320: data = 8'hfe;
      17'd44321: data = 8'hfd;
      17'd44322: data = 8'hfd;
      17'd44323: data = 8'hfd;
      17'd44324: data = 8'hfd;
      17'd44325: data = 8'hfe;
      17'd44326: data = 8'hfd;
      17'd44327: data = 8'hfe;
      17'd44328: data = 8'hfe;
      17'd44329: data = 8'h00;
      17'd44330: data = 8'h00;
      17'd44331: data = 8'h00;
      17'd44332: data = 8'h00;
      17'd44333: data = 8'h01;
      17'd44334: data = 8'h00;
      17'd44335: data = 8'h00;
      17'd44336: data = 8'h01;
      17'd44337: data = 8'h00;
      17'd44338: data = 8'hfe;
      17'd44339: data = 8'h00;
      17'd44340: data = 8'h00;
      17'd44341: data = 8'h00;
      17'd44342: data = 8'h01;
      17'd44343: data = 8'h01;
      17'd44344: data = 8'h00;
      17'd44345: data = 8'h00;
      17'd44346: data = 8'h01;
      17'd44347: data = 8'h01;
      17'd44348: data = 8'h00;
      17'd44349: data = 8'h01;
      17'd44350: data = 8'h02;
      17'd44351: data = 8'h00;
      17'd44352: data = 8'h00;
      17'd44353: data = 8'h01;
      17'd44354: data = 8'h00;
      17'd44355: data = 8'hfe;
      17'd44356: data = 8'h00;
      17'd44357: data = 8'h00;
      17'd44358: data = 8'h00;
      17'd44359: data = 8'h01;
      17'd44360: data = 8'hfe;
      17'd44361: data = 8'h00;
      17'd44362: data = 8'h01;
      17'd44363: data = 8'h01;
      17'd44364: data = 8'hfe;
      17'd44365: data = 8'hfe;
      17'd44366: data = 8'h00;
      17'd44367: data = 8'h00;
      17'd44368: data = 8'h00;
      17'd44369: data = 8'h00;
      17'd44370: data = 8'hfe;
      17'd44371: data = 8'h00;
      17'd44372: data = 8'h02;
      17'd44373: data = 8'h01;
      17'd44374: data = 8'h01;
      17'd44375: data = 8'h02;
      17'd44376: data = 8'h01;
      17'd44377: data = 8'h01;
      17'd44378: data = 8'h04;
      17'd44379: data = 8'h01;
      17'd44380: data = 8'hfe;
      17'd44381: data = 8'h00;
      17'd44382: data = 8'h00;
      17'd44383: data = 8'h00;
      17'd44384: data = 8'h00;
      17'd44385: data = 8'h00;
      17'd44386: data = 8'hfe;
      17'd44387: data = 8'h01;
      17'd44388: data = 8'h04;
      17'd44389: data = 8'h01;
      17'd44390: data = 8'h00;
      17'd44391: data = 8'h01;
      17'd44392: data = 8'h04;
      17'd44393: data = 8'h02;
      17'd44394: data = 8'h00;
      17'd44395: data = 8'h02;
      17'd44396: data = 8'h01;
      17'd44397: data = 8'h04;
      17'd44398: data = 8'h02;
      17'd44399: data = 8'h00;
      17'd44400: data = 8'h00;
      17'd44401: data = 8'hfe;
      17'd44402: data = 8'h01;
      17'd44403: data = 8'h02;
      17'd44404: data = 8'h00;
      17'd44405: data = 8'h00;
      17'd44406: data = 8'h01;
      17'd44407: data = 8'h02;
      17'd44408: data = 8'h02;
      17'd44409: data = 8'h01;
      17'd44410: data = 8'h00;
      17'd44411: data = 8'h00;
      17'd44412: data = 8'h01;
      17'd44413: data = 8'h00;
      17'd44414: data = 8'hfd;
      17'd44415: data = 8'hfd;
      17'd44416: data = 8'hfd;
      17'd44417: data = 8'h00;
      17'd44418: data = 8'h00;
      17'd44419: data = 8'hfd;
      17'd44420: data = 8'hfd;
      17'd44421: data = 8'hfe;
      17'd44422: data = 8'h00;
      17'd44423: data = 8'h00;
      17'd44424: data = 8'hfd;
      17'd44425: data = 8'hfd;
      17'd44426: data = 8'h00;
      17'd44427: data = 8'h00;
      17'd44428: data = 8'hfe;
      17'd44429: data = 8'hfd;
      17'd44430: data = 8'hfe;
      17'd44431: data = 8'h00;
      17'd44432: data = 8'hfd;
      17'd44433: data = 8'hfe;
      17'd44434: data = 8'hfe;
      17'd44435: data = 8'hfd;
      17'd44436: data = 8'h00;
      17'd44437: data = 8'h00;
      17'd44438: data = 8'hfe;
      17'd44439: data = 8'h01;
      17'd44440: data = 8'h01;
      17'd44441: data = 8'h00;
      17'd44442: data = 8'h00;
      17'd44443: data = 8'h00;
      17'd44444: data = 8'h00;
      17'd44445: data = 8'h00;
      17'd44446: data = 8'h02;
      17'd44447: data = 8'h01;
      17'd44448: data = 8'h00;
      17'd44449: data = 8'h00;
      17'd44450: data = 8'h01;
      17'd44451: data = 8'h00;
      17'd44452: data = 8'hfe;
      17'd44453: data = 8'hfe;
      17'd44454: data = 8'h00;
      17'd44455: data = 8'h01;
      17'd44456: data = 8'h01;
      17'd44457: data = 8'hfe;
      17'd44458: data = 8'hfe;
      17'd44459: data = 8'hfe;
      17'd44460: data = 8'h00;
      17'd44461: data = 8'h01;
      17'd44462: data = 8'hfd;
      17'd44463: data = 8'hfe;
      17'd44464: data = 8'h00;
      17'd44465: data = 8'hfe;
      17'd44466: data = 8'h00;
      17'd44467: data = 8'h00;
      17'd44468: data = 8'hfe;
      17'd44469: data = 8'h00;
      17'd44470: data = 8'h00;
      17'd44471: data = 8'hfe;
      17'd44472: data = 8'hfe;
      17'd44473: data = 8'hfe;
      17'd44474: data = 8'hfd;
      17'd44475: data = 8'hfe;
      17'd44476: data = 8'hfe;
      17'd44477: data = 8'hfa;
      17'd44478: data = 8'hfd;
      17'd44479: data = 8'hfe;
      17'd44480: data = 8'hfe;
      17'd44481: data = 8'hfc;
      17'd44482: data = 8'hfd;
      17'd44483: data = 8'hfd;
      17'd44484: data = 8'hfe;
      17'd44485: data = 8'h00;
      17'd44486: data = 8'hfe;
      17'd44487: data = 8'hfe;
      17'd44488: data = 8'h00;
      17'd44489: data = 8'h00;
      17'd44490: data = 8'hfe;
      17'd44491: data = 8'h00;
      17'd44492: data = 8'hfd;
      17'd44493: data = 8'hfe;
      17'd44494: data = 8'h02;
      17'd44495: data = 8'h00;
      17'd44496: data = 8'h00;
      17'd44497: data = 8'h00;
      17'd44498: data = 8'h00;
      17'd44499: data = 8'h01;
      17'd44500: data = 8'h01;
      17'd44501: data = 8'h00;
      17'd44502: data = 8'h00;
      17'd44503: data = 8'h01;
      17'd44504: data = 8'h01;
      17'd44505: data = 8'h00;
      17'd44506: data = 8'hfe;
      17'd44507: data = 8'hfd;
      17'd44508: data = 8'hfe;
      17'd44509: data = 8'h00;
      17'd44510: data = 8'hfd;
      17'd44511: data = 8'hfd;
      17'd44512: data = 8'hfd;
      17'd44513: data = 8'hfd;
      17'd44514: data = 8'hfd;
      17'd44515: data = 8'hfd;
      17'd44516: data = 8'hfa;
      17'd44517: data = 8'hfa;
      17'd44518: data = 8'hfd;
      17'd44519: data = 8'hfe;
      17'd44520: data = 8'hfe;
      17'd44521: data = 8'hfd;
      17'd44522: data = 8'hfd;
      17'd44523: data = 8'h00;
      17'd44524: data = 8'hfe;
      17'd44525: data = 8'hfd;
      17'd44526: data = 8'hfd;
      17'd44527: data = 8'hfd;
      17'd44528: data = 8'hfd;
      17'd44529: data = 8'hfd;
      17'd44530: data = 8'hfe;
      17'd44531: data = 8'hfe;
      17'd44532: data = 8'hfd;
      17'd44533: data = 8'h00;
      17'd44534: data = 8'h00;
      17'd44535: data = 8'h00;
      17'd44536: data = 8'hfe;
      17'd44537: data = 8'hfe;
      17'd44538: data = 8'hfe;
      17'd44539: data = 8'h01;
      17'd44540: data = 8'hfe;
      17'd44541: data = 8'hfe;
      17'd44542: data = 8'h00;
      17'd44543: data = 8'h00;
      17'd44544: data = 8'hfe;
      17'd44545: data = 8'hfd;
      17'd44546: data = 8'hfe;
      17'd44547: data = 8'hfd;
      17'd44548: data = 8'hfe;
      17'd44549: data = 8'h00;
      17'd44550: data = 8'hfe;
      17'd44551: data = 8'hfc;
      17'd44552: data = 8'hfe;
      17'd44553: data = 8'h01;
      17'd44554: data = 8'hfe;
      17'd44555: data = 8'hfd;
      17'd44556: data = 8'hfd;
      17'd44557: data = 8'hfd;
      17'd44558: data = 8'hfd;
      17'd44559: data = 8'hfd;
      17'd44560: data = 8'hfe;
      17'd44561: data = 8'hfd;
      17'd44562: data = 8'hfd;
      17'd44563: data = 8'hfe;
      17'd44564: data = 8'hfe;
      17'd44565: data = 8'hfe;
      17'd44566: data = 8'hfe;
      17'd44567: data = 8'h00;
      17'd44568: data = 8'h01;
      17'd44569: data = 8'h00;
      17'd44570: data = 8'hfd;
      17'd44571: data = 8'hfe;
      17'd44572: data = 8'h00;
      17'd44573: data = 8'h00;
      17'd44574: data = 8'hfd;
      17'd44575: data = 8'hfe;
      17'd44576: data = 8'h00;
      17'd44577: data = 8'h00;
      17'd44578: data = 8'h01;
      17'd44579: data = 8'hfe;
      17'd44580: data = 8'hfe;
      17'd44581: data = 8'h00;
      17'd44582: data = 8'h01;
      17'd44583: data = 8'h00;
      17'd44584: data = 8'hfe;
      17'd44585: data = 8'h00;
      17'd44586: data = 8'hfe;
      17'd44587: data = 8'hfe;
      17'd44588: data = 8'h00;
      17'd44589: data = 8'hfe;
      17'd44590: data = 8'hfe;
      17'd44591: data = 8'hfd;
      17'd44592: data = 8'h00;
      17'd44593: data = 8'h00;
      17'd44594: data = 8'hfe;
      17'd44595: data = 8'hfe;
      17'd44596: data = 8'hfe;
      17'd44597: data = 8'h01;
      17'd44598: data = 8'h00;
      17'd44599: data = 8'hfe;
      17'd44600: data = 8'hfe;
      17'd44601: data = 8'hfd;
      17'd44602: data = 8'h00;
      17'd44603: data = 8'hfe;
      17'd44604: data = 8'hfc;
      17'd44605: data = 8'hfc;
      17'd44606: data = 8'hfd;
      17'd44607: data = 8'hfe;
      17'd44608: data = 8'h00;
      17'd44609: data = 8'hfe;
      17'd44610: data = 8'hfc;
      17'd44611: data = 8'hfd;
      17'd44612: data = 8'h01;
      17'd44613: data = 8'h00;
      17'd44614: data = 8'hfe;
      17'd44615: data = 8'h00;
      17'd44616: data = 8'h00;
      17'd44617: data = 8'hfe;
      17'd44618: data = 8'h01;
      17'd44619: data = 8'h00;
      17'd44620: data = 8'hfe;
      17'd44621: data = 8'hfd;
      17'd44622: data = 8'hfd;
      17'd44623: data = 8'hfe;
      17'd44624: data = 8'h00;
      17'd44625: data = 8'hfe;
      17'd44626: data = 8'hfe;
      17'd44627: data = 8'hfe;
      17'd44628: data = 8'h00;
      17'd44629: data = 8'h01;
      17'd44630: data = 8'hfe;
      17'd44631: data = 8'h00;
      17'd44632: data = 8'h02;
      17'd44633: data = 8'h01;
      17'd44634: data = 8'h00;
      17'd44635: data = 8'h01;
      17'd44636: data = 8'h02;
      17'd44637: data = 8'h01;
      17'd44638: data = 8'h02;
      17'd44639: data = 8'h00;
      17'd44640: data = 8'h00;
      17'd44641: data = 8'h00;
      17'd44642: data = 8'h01;
      17'd44643: data = 8'h00;
      17'd44644: data = 8'hfe;
      17'd44645: data = 8'h02;
      17'd44646: data = 8'h01;
      17'd44647: data = 8'h01;
      17'd44648: data = 8'h01;
      17'd44649: data = 8'hfd;
      17'd44650: data = 8'h00;
      17'd44651: data = 8'h02;
      17'd44652: data = 8'hfe;
      17'd44653: data = 8'hfe;
      17'd44654: data = 8'h00;
      17'd44655: data = 8'h00;
      17'd44656: data = 8'h01;
      17'd44657: data = 8'h02;
      17'd44658: data = 8'h01;
      17'd44659: data = 8'h01;
      17'd44660: data = 8'h01;
      17'd44661: data = 8'h02;
      17'd44662: data = 8'h04;
      17'd44663: data = 8'h01;
      17'd44664: data = 8'h02;
      17'd44665: data = 8'h01;
      17'd44666: data = 8'h01;
      17'd44667: data = 8'h01;
      17'd44668: data = 8'hfd;
      17'd44669: data = 8'hfd;
      17'd44670: data = 8'hfe;
      17'd44671: data = 8'h01;
      17'd44672: data = 8'h00;
      17'd44673: data = 8'hfd;
      17'd44674: data = 8'h00;
      17'd44675: data = 8'h01;
      17'd44676: data = 8'h00;
      17'd44677: data = 8'h00;
      17'd44678: data = 8'hfe;
      17'd44679: data = 8'hfe;
      17'd44680: data = 8'h00;
      17'd44681: data = 8'h00;
      17'd44682: data = 8'hfd;
      17'd44683: data = 8'hfc;
      17'd44684: data = 8'hfd;
      17'd44685: data = 8'hfd;
      17'd44686: data = 8'hfd;
      17'd44687: data = 8'hfd;
      17'd44688: data = 8'hfd;
      17'd44689: data = 8'hfc;
      17'd44690: data = 8'hfe;
      17'd44691: data = 8'hfe;
      17'd44692: data = 8'h00;
      17'd44693: data = 8'hfe;
      17'd44694: data = 8'hfe;
      17'd44695: data = 8'h00;
      17'd44696: data = 8'hfe;
      17'd44697: data = 8'hfe;
      17'd44698: data = 8'hfd;
      17'd44699: data = 8'hfd;
      17'd44700: data = 8'hfc;
      17'd44701: data = 8'hfc;
      17'd44702: data = 8'hfd;
      17'd44703: data = 8'hfe;
      17'd44704: data = 8'hfd;
      17'd44705: data = 8'hfe;
      17'd44706: data = 8'hfe;
      17'd44707: data = 8'h00;
      17'd44708: data = 8'h00;
      17'd44709: data = 8'h00;
      17'd44710: data = 8'h00;
      17'd44711: data = 8'hfe;
      17'd44712: data = 8'hfe;
      17'd44713: data = 8'h00;
      17'd44714: data = 8'h00;
      17'd44715: data = 8'h00;
      17'd44716: data = 8'hfe;
      17'd44717: data = 8'hfe;
      17'd44718: data = 8'h00;
      17'd44719: data = 8'h00;
      17'd44720: data = 8'hfe;
      17'd44721: data = 8'h00;
      17'd44722: data = 8'h01;
      17'd44723: data = 8'h00;
      17'd44724: data = 8'h01;
      17'd44725: data = 8'h00;
      17'd44726: data = 8'hfe;
      17'd44727: data = 8'hfe;
      17'd44728: data = 8'h00;
      17'd44729: data = 8'h00;
      17'd44730: data = 8'hfe;
      17'd44731: data = 8'hfe;
      17'd44732: data = 8'hfe;
      17'd44733: data = 8'hfe;
      17'd44734: data = 8'h00;
      17'd44735: data = 8'h01;
      17'd44736: data = 8'h00;
      17'd44737: data = 8'hfd;
      17'd44738: data = 8'h00;
      17'd44739: data = 8'h02;
      17'd44740: data = 8'h00;
      17'd44741: data = 8'h00;
      17'd44742: data = 8'h00;
      17'd44743: data = 8'hfe;
      17'd44744: data = 8'hfe;
      17'd44745: data = 8'hfe;
      17'd44746: data = 8'hfe;
      17'd44747: data = 8'hfd;
      17'd44748: data = 8'hfe;
      17'd44749: data = 8'hfe;
      17'd44750: data = 8'h00;
      17'd44751: data = 8'hfd;
      17'd44752: data = 8'hfd;
      17'd44753: data = 8'hfe;
      17'd44754: data = 8'h00;
      17'd44755: data = 8'hfe;
      17'd44756: data = 8'h00;
      17'd44757: data = 8'hfe;
      17'd44758: data = 8'hfd;
      17'd44759: data = 8'hfe;
      17'd44760: data = 8'h01;
      17'd44761: data = 8'h06;
      17'd44762: data = 8'h05;
      17'd44763: data = 8'hfc;
      17'd44764: data = 8'hf9;
      17'd44765: data = 8'hfe;
      17'd44766: data = 8'h00;
      17'd44767: data = 8'h01;
      17'd44768: data = 8'hfe;
      17'd44769: data = 8'hfd;
      17'd44770: data = 8'h02;
      17'd44771: data = 8'h05;
      17'd44772: data = 8'hfe;
      17'd44773: data = 8'hfc;
      17'd44774: data = 8'h01;
      17'd44775: data = 8'h05;
      17'd44776: data = 8'h02;
      17'd44777: data = 8'hfd;
      17'd44778: data = 8'hfa;
      17'd44779: data = 8'hfd;
      17'd44780: data = 8'h04;
      17'd44781: data = 8'h05;
      17'd44782: data = 8'hfc;
      17'd44783: data = 8'hf9;
      17'd44784: data = 8'hfc;
      17'd44785: data = 8'h00;
      17'd44786: data = 8'hfd;
      17'd44787: data = 8'hfa;
      17'd44788: data = 8'hfd;
      17'd44789: data = 8'hfe;
      17'd44790: data = 8'h01;
      17'd44791: data = 8'h00;
      17'd44792: data = 8'hfd;
      17'd44793: data = 8'hfe;
      17'd44794: data = 8'h02;
      17'd44795: data = 8'h02;
      17'd44796: data = 8'hfe;
      17'd44797: data = 8'hfc;
      17'd44798: data = 8'hfa;
      17'd44799: data = 8'h00;
      17'd44800: data = 8'h00;
      17'd44801: data = 8'hfe;
      17'd44802: data = 8'hfc;
      17'd44803: data = 8'hfe;
      17'd44804: data = 8'h04;
      17'd44805: data = 8'h01;
      17'd44806: data = 8'hfe;
      17'd44807: data = 8'hfe;
      17'd44808: data = 8'h02;
      17'd44809: data = 8'h00;
      17'd44810: data = 8'hfd;
      17'd44811: data = 8'hfc;
      17'd44812: data = 8'hfc;
      17'd44813: data = 8'h00;
      17'd44814: data = 8'h01;
      17'd44815: data = 8'h00;
      17'd44816: data = 8'h00;
      17'd44817: data = 8'hfe;
      17'd44818: data = 8'h00;
      17'd44819: data = 8'h02;
      17'd44820: data = 8'h02;
      17'd44821: data = 8'h00;
      17'd44822: data = 8'h00;
      17'd44823: data = 8'h01;
      17'd44824: data = 8'h02;
      17'd44825: data = 8'h02;
      17'd44826: data = 8'h00;
      17'd44827: data = 8'hfe;
      17'd44828: data = 8'h00;
      17'd44829: data = 8'h00;
      17'd44830: data = 8'h00;
      17'd44831: data = 8'hfe;
      17'd44832: data = 8'h00;
      17'd44833: data = 8'h00;
      17'd44834: data = 8'h00;
      17'd44835: data = 8'h02;
      17'd44836: data = 8'h02;
      17'd44837: data = 8'h00;
      17'd44838: data = 8'h00;
      17'd44839: data = 8'h01;
      17'd44840: data = 8'h00;
      17'd44841: data = 8'h00;
      17'd44842: data = 8'h00;
      17'd44843: data = 8'hfd;
      17'd44844: data = 8'hfd;
      17'd44845: data = 8'hfd;
      17'd44846: data = 8'hfc;
      17'd44847: data = 8'hfe;
      17'd44848: data = 8'hfd;
      17'd44849: data = 8'h00;
      17'd44850: data = 8'h00;
      17'd44851: data = 8'h00;
      17'd44852: data = 8'h02;
      17'd44853: data = 8'h00;
      17'd44854: data = 8'h00;
      17'd44855: data = 8'h00;
      17'd44856: data = 8'hfe;
      17'd44857: data = 8'h00;
      17'd44858: data = 8'h00;
      17'd44859: data = 8'h01;
      17'd44860: data = 8'h01;
      17'd44861: data = 8'h00;
      17'd44862: data = 8'h00;
      17'd44863: data = 8'h01;
      17'd44864: data = 8'h01;
      17'd44865: data = 8'h02;
      17'd44866: data = 8'h00;
      17'd44867: data = 8'h01;
      17'd44868: data = 8'h01;
      17'd44869: data = 8'h01;
      17'd44870: data = 8'h02;
      17'd44871: data = 8'hfe;
      17'd44872: data = 8'hfe;
      17'd44873: data = 8'h00;
      17'd44874: data = 8'h00;
      17'd44875: data = 8'h00;
      17'd44876: data = 8'h00;
      17'd44877: data = 8'h01;
      17'd44878: data = 8'h00;
      17'd44879: data = 8'hfe;
      17'd44880: data = 8'h02;
      17'd44881: data = 8'h02;
      17'd44882: data = 8'hfe;
      17'd44883: data = 8'h00;
      17'd44884: data = 8'h00;
      17'd44885: data = 8'h01;
      17'd44886: data = 8'h00;
      17'd44887: data = 8'hfe;
      17'd44888: data = 8'hfd;
      17'd44889: data = 8'hfd;
      17'd44890: data = 8'h00;
      17'd44891: data = 8'hfe;
      17'd44892: data = 8'hfe;
      17'd44893: data = 8'hfe;
      17'd44894: data = 8'hfe;
      17'd44895: data = 8'hfe;
      17'd44896: data = 8'h00;
      17'd44897: data = 8'h01;
      17'd44898: data = 8'h01;
      17'd44899: data = 8'h00;
      17'd44900: data = 8'hfe;
      17'd44901: data = 8'hfc;
      17'd44902: data = 8'hfd;
      17'd44903: data = 8'hfd;
      17'd44904: data = 8'hfd;
      17'd44905: data = 8'hfd;
      17'd44906: data = 8'hfc;
      17'd44907: data = 8'hfd;
      17'd44908: data = 8'h00;
      17'd44909: data = 8'hfe;
      17'd44910: data = 8'hfe;
      17'd44911: data = 8'hfd;
      17'd44912: data = 8'hfe;
      17'd44913: data = 8'h00;
      17'd44914: data = 8'h00;
      17'd44915: data = 8'hfe;
      17'd44916: data = 8'hfc;
      17'd44917: data = 8'hfe;
      17'd44918: data = 8'hfe;
      17'd44919: data = 8'hfe;
      17'd44920: data = 8'hfd;
      17'd44921: data = 8'hfe;
      17'd44922: data = 8'h00;
      17'd44923: data = 8'h00;
      17'd44924: data = 8'h01;
      17'd44925: data = 8'h01;
      17'd44926: data = 8'h00;
      17'd44927: data = 8'h00;
      17'd44928: data = 8'h00;
      17'd44929: data = 8'h00;
      17'd44930: data = 8'hfe;
      17'd44931: data = 8'h00;
      17'd44932: data = 8'hfe;
      17'd44933: data = 8'hfe;
      17'd44934: data = 8'hfe;
      17'd44935: data = 8'hfe;
      17'd44936: data = 8'hfe;
      17'd44937: data = 8'h00;
      17'd44938: data = 8'h01;
      17'd44939: data = 8'h01;
      17'd44940: data = 8'h01;
      17'd44941: data = 8'h00;
      17'd44942: data = 8'h01;
      17'd44943: data = 8'h02;
      17'd44944: data = 8'h00;
      17'd44945: data = 8'hfd;
      17'd44946: data = 8'hfd;
      17'd44947: data = 8'hfe;
      17'd44948: data = 8'h00;
      17'd44949: data = 8'hfe;
      17'd44950: data = 8'hfe;
      17'd44951: data = 8'hfc;
      17'd44952: data = 8'hfe;
      17'd44953: data = 8'h01;
      17'd44954: data = 8'h00;
      17'd44955: data = 8'hfe;
      17'd44956: data = 8'h00;
      17'd44957: data = 8'h01;
      17'd44958: data = 8'h00;
      17'd44959: data = 8'h00;
      17'd44960: data = 8'hfc;
      17'd44961: data = 8'hfd;
      17'd44962: data = 8'hfd;
      17'd44963: data = 8'hfd;
      17'd44964: data = 8'hfd;
      17'd44965: data = 8'hfd;
      17'd44966: data = 8'hfe;
      17'd44967: data = 8'hfe;
      17'd44968: data = 8'hfe;
      17'd44969: data = 8'hfe;
      17'd44970: data = 8'h00;
      17'd44971: data = 8'h02;
      17'd44972: data = 8'h01;
      17'd44973: data = 8'h00;
      17'd44974: data = 8'hfe;
      17'd44975: data = 8'hfe;
      17'd44976: data = 8'h01;
      17'd44977: data = 8'h00;
      17'd44978: data = 8'hfe;
      17'd44979: data = 8'hfc;
      17'd44980: data = 8'hfe;
      17'd44981: data = 8'h00;
      17'd44982: data = 8'h00;
      17'd44983: data = 8'hfe;
      17'd44984: data = 8'hfd;
      17'd44985: data = 8'hfe;
      17'd44986: data = 8'h00;
      17'd44987: data = 8'h01;
      17'd44988: data = 8'hfd;
      17'd44989: data = 8'hfc;
      17'd44990: data = 8'hfe;
      17'd44991: data = 8'h00;
      17'd44992: data = 8'hfe;
      17'd44993: data = 8'hfe;
      17'd44994: data = 8'hfd;
      17'd44995: data = 8'hfe;
      17'd44996: data = 8'h01;
      17'd44997: data = 8'h01;
      17'd44998: data = 8'hfe;
      17'd44999: data = 8'h00;
      17'd45000: data = 8'h04;
      17'd45001: data = 8'h02;
      17'd45002: data = 8'h01;
      17'd45003: data = 8'h00;
      17'd45004: data = 8'h01;
      17'd45005: data = 8'h04;
      17'd45006: data = 8'h01;
      17'd45007: data = 8'h00;
      17'd45008: data = 8'hfe;
      17'd45009: data = 8'hfe;
      17'd45010: data = 8'h01;
      17'd45011: data = 8'h00;
      17'd45012: data = 8'hfd;
      17'd45013: data = 8'hfe;
      17'd45014: data = 8'h00;
      17'd45015: data = 8'h01;
      17'd45016: data = 8'h00;
      17'd45017: data = 8'h00;
      17'd45018: data = 8'h00;
      17'd45019: data = 8'h01;
      17'd45020: data = 8'h02;
      17'd45021: data = 8'h00;
      17'd45022: data = 8'h00;
      17'd45023: data = 8'h00;
      17'd45024: data = 8'h00;
      17'd45025: data = 8'h01;
      17'd45026: data = 8'h00;
      17'd45027: data = 8'hfc;
      17'd45028: data = 8'hfe;
      17'd45029: data = 8'h06;
      17'd45030: data = 8'hfe;
      17'd45031: data = 8'hf6;
      17'd45032: data = 8'hfe;
      17'd45033: data = 8'hfe;
      17'd45034: data = 8'hfe;
      17'd45035: data = 8'hfd;
      17'd45036: data = 8'hf9;
      17'd45037: data = 8'h01;
      17'd45038: data = 8'h05;
      17'd45039: data = 8'hfd;
      17'd45040: data = 8'hf9;
      17'd45041: data = 8'hfe;
      17'd45042: data = 8'h04;
      17'd45043: data = 8'hfe;
      17'd45044: data = 8'hfa;
      17'd45045: data = 8'hfa;
      17'd45046: data = 8'hfe;
      17'd45047: data = 8'hfe;
      17'd45048: data = 8'hfe;
      17'd45049: data = 8'hfd;
      17'd45050: data = 8'hfc;
      17'd45051: data = 8'h04;
      17'd45052: data = 8'h01;
      17'd45053: data = 8'hfc;
      17'd45054: data = 8'hfe;
      17'd45055: data = 8'h02;
      17'd45056: data = 8'h04;
      17'd45057: data = 8'hfe;
      17'd45058: data = 8'hfd;
      17'd45059: data = 8'h01;
      17'd45060: data = 8'h00;
      17'd45061: data = 8'h00;
      17'd45062: data = 8'h00;
      17'd45063: data = 8'h01;
      17'd45064: data = 8'h00;
      17'd45065: data = 8'hfe;
      17'd45066: data = 8'hfe;
      17'd45067: data = 8'h02;
      17'd45068: data = 8'h00;
      17'd45069: data = 8'hfd;
      17'd45070: data = 8'hfd;
      17'd45071: data = 8'h00;
      17'd45072: data = 8'h04;
      17'd45073: data = 8'hfe;
      17'd45074: data = 8'hfc;
      17'd45075: data = 8'h00;
      17'd45076: data = 8'h04;
      17'd45077: data = 8'h01;
      17'd45078: data = 8'hfd;
      17'd45079: data = 8'hfe;
      17'd45080: data = 8'h00;
      17'd45081: data = 8'h01;
      17'd45082: data = 8'hfd;
      17'd45083: data = 8'hfa;
      17'd45084: data = 8'hfd;
      17'd45085: data = 8'h01;
      17'd45086: data = 8'h00;
      17'd45087: data = 8'hfa;
      17'd45088: data = 8'h00;
      17'd45089: data = 8'h02;
      17'd45090: data = 8'hfe;
      17'd45091: data = 8'hfd;
      17'd45092: data = 8'hfd;
      17'd45093: data = 8'h00;
      17'd45094: data = 8'h00;
      17'd45095: data = 8'hfd;
      17'd45096: data = 8'hfe;
      17'd45097: data = 8'hfe;
      17'd45098: data = 8'h01;
      17'd45099: data = 8'h01;
      17'd45100: data = 8'hfe;
      17'd45101: data = 8'hfe;
      17'd45102: data = 8'h01;
      17'd45103: data = 8'h00;
      17'd45104: data = 8'h00;
      17'd45105: data = 8'h00;
      17'd45106: data = 8'hfd;
      17'd45107: data = 8'hfd;
      17'd45108: data = 8'hfe;
      17'd45109: data = 8'h00;
      17'd45110: data = 8'h00;
      17'd45111: data = 8'hfe;
      17'd45112: data = 8'hfe;
      17'd45113: data = 8'hfe;
      17'd45114: data = 8'hfe;
      17'd45115: data = 8'h00;
      17'd45116: data = 8'hfe;
      17'd45117: data = 8'hfe;
      17'd45118: data = 8'h00;
      17'd45119: data = 8'h00;
      17'd45120: data = 8'h01;
      17'd45121: data = 8'h00;
      17'd45122: data = 8'hfe;
      17'd45123: data = 8'h00;
      17'd45124: data = 8'h00;
      17'd45125: data = 8'h00;
      17'd45126: data = 8'h00;
      17'd45127: data = 8'hfe;
      17'd45128: data = 8'h00;
      17'd45129: data = 8'h00;
      17'd45130: data = 8'h01;
      17'd45131: data = 8'h00;
      17'd45132: data = 8'h00;
      17'd45133: data = 8'h01;
      17'd45134: data = 8'h01;
      17'd45135: data = 8'h01;
      17'd45136: data = 8'h02;
      17'd45137: data = 8'h02;
      17'd45138: data = 8'h00;
      17'd45139: data = 8'h00;
      17'd45140: data = 8'h00;
      17'd45141: data = 8'hfe;
      17'd45142: data = 8'hfe;
      17'd45143: data = 8'hfd;
      17'd45144: data = 8'hfe;
      17'd45145: data = 8'h00;
      17'd45146: data = 8'h01;
      17'd45147: data = 8'h00;
      17'd45148: data = 8'h00;
      17'd45149: data = 8'h01;
      17'd45150: data = 8'h01;
      17'd45151: data = 8'h00;
      17'd45152: data = 8'h01;
      17'd45153: data = 8'h01;
      17'd45154: data = 8'h01;
      17'd45155: data = 8'h01;
      17'd45156: data = 8'h00;
      17'd45157: data = 8'hfe;
      17'd45158: data = 8'hfd;
      17'd45159: data = 8'h00;
      17'd45160: data = 8'h00;
      17'd45161: data = 8'h00;
      17'd45162: data = 8'h00;
      17'd45163: data = 8'h01;
      17'd45164: data = 8'h01;
      17'd45165: data = 8'h00;
      17'd45166: data = 8'h01;
      17'd45167: data = 8'h00;
      17'd45168: data = 8'hfe;
      17'd45169: data = 8'hfe;
      17'd45170: data = 8'h00;
      17'd45171: data = 8'hfe;
      17'd45172: data = 8'hfe;
      17'd45173: data = 8'hfe;
      17'd45174: data = 8'hfe;
      17'd45175: data = 8'h00;
      17'd45176: data = 8'h01;
      17'd45177: data = 8'h01;
      17'd45178: data = 8'h01;
      17'd45179: data = 8'h01;
      17'd45180: data = 8'h01;
      17'd45181: data = 8'h01;
      17'd45182: data = 8'h02;
      17'd45183: data = 8'h01;
      17'd45184: data = 8'h02;
      17'd45185: data = 8'h02;
      17'd45186: data = 8'h01;
      17'd45187: data = 8'h02;
      17'd45188: data = 8'h02;
      17'd45189: data = 8'h01;
      17'd45190: data = 8'h02;
      17'd45191: data = 8'h01;
      17'd45192: data = 8'h01;
      17'd45193: data = 8'h02;
      17'd45194: data = 8'h02;
      17'd45195: data = 8'h02;
      17'd45196: data = 8'h02;
      17'd45197: data = 8'h02;
      17'd45198: data = 8'h01;
      17'd45199: data = 8'h02;
      17'd45200: data = 8'h02;
      17'd45201: data = 8'h01;
      17'd45202: data = 8'hfe;
      17'd45203: data = 8'h00;
      17'd45204: data = 8'h00;
      17'd45205: data = 8'hfe;
      17'd45206: data = 8'hfe;
      17'd45207: data = 8'hfe;
      17'd45208: data = 8'hfe;
      17'd45209: data = 8'h00;
      17'd45210: data = 8'h00;
      17'd45211: data = 8'hfe;
      17'd45212: data = 8'hfe;
      17'd45213: data = 8'h00;
      17'd45214: data = 8'h01;
      17'd45215: data = 8'h01;
      17'd45216: data = 8'h00;
      17'd45217: data = 8'hfe;
      17'd45218: data = 8'h00;
      17'd45219: data = 8'h01;
      17'd45220: data = 8'h01;
      17'd45221: data = 8'hfe;
      17'd45222: data = 8'hfe;
      17'd45223: data = 8'hfe;
      17'd45224: data = 8'h01;
      17'd45225: data = 8'h01;
      17'd45226: data = 8'hfd;
      17'd45227: data = 8'hfd;
      17'd45228: data = 8'h00;
      17'd45229: data = 8'hfe;
      17'd45230: data = 8'hfe;
      17'd45231: data = 8'hfe;
      17'd45232: data = 8'hfe;
      17'd45233: data = 8'hfe;
      17'd45234: data = 8'h02;
      17'd45235: data = 8'h01;
      17'd45236: data = 8'h00;
      17'd45237: data = 8'h01;
      17'd45238: data = 8'h01;
      17'd45239: data = 8'h00;
      17'd45240: data = 8'h00;
      17'd45241: data = 8'hfe;
      17'd45242: data = 8'h00;
      17'd45243: data = 8'h01;
      17'd45244: data = 8'hfe;
      17'd45245: data = 8'h00;
      17'd45246: data = 8'h00;
      17'd45247: data = 8'h00;
      17'd45248: data = 8'h02;
      17'd45249: data = 8'h01;
      17'd45250: data = 8'h00;
      17'd45251: data = 8'h01;
      17'd45252: data = 8'h01;
      17'd45253: data = 8'h02;
      17'd45254: data = 8'h01;
      17'd45255: data = 8'h00;
      17'd45256: data = 8'hfd;
      17'd45257: data = 8'h00;
      17'd45258: data = 8'h00;
      17'd45259: data = 8'hfe;
      17'd45260: data = 8'hfe;
      17'd45261: data = 8'h00;
      17'd45262: data = 8'h01;
      17'd45263: data = 8'h02;
      17'd45264: data = 8'h01;
      17'd45265: data = 8'h01;
      17'd45266: data = 8'h01;
      17'd45267: data = 8'h00;
      17'd45268: data = 8'h00;
      17'd45269: data = 8'h00;
      17'd45270: data = 8'hfe;
      17'd45271: data = 8'hfd;
      17'd45272: data = 8'hfe;
      17'd45273: data = 8'hfe;
      17'd45274: data = 8'hfe;
      17'd45275: data = 8'hfe;
      17'd45276: data = 8'hfe;
      17'd45277: data = 8'h01;
      17'd45278: data = 8'h02;
      17'd45279: data = 8'h01;
      17'd45280: data = 8'h01;
      17'd45281: data = 8'h02;
      17'd45282: data = 8'h02;
      17'd45283: data = 8'h00;
      17'd45284: data = 8'hfe;
      17'd45285: data = 8'hfe;
      17'd45286: data = 8'hfd;
      17'd45287: data = 8'hfd;
      17'd45288: data = 8'hfd;
      17'd45289: data = 8'hfd;
      17'd45290: data = 8'hfe;
      17'd45291: data = 8'h01;
      17'd45292: data = 8'h01;
      17'd45293: data = 8'h00;
      17'd45294: data = 8'h00;
      17'd45295: data = 8'h01;
      17'd45296: data = 8'h01;
      17'd45297: data = 8'h00;
      17'd45298: data = 8'h00;
      17'd45299: data = 8'h00;
      17'd45300: data = 8'hfe;
      17'd45301: data = 8'h00;
      17'd45302: data = 8'hfd;
      17'd45303: data = 8'hfe;
      17'd45304: data = 8'h00;
      17'd45305: data = 8'hfe;
      17'd45306: data = 8'hfe;
      17'd45307: data = 8'h00;
      17'd45308: data = 8'h00;
      17'd45309: data = 8'h01;
      17'd45310: data = 8'h00;
      17'd45311: data = 8'h00;
      17'd45312: data = 8'h00;
      17'd45313: data = 8'h01;
      17'd45314: data = 8'h01;
      17'd45315: data = 8'h01;
      17'd45316: data = 8'h01;
      17'd45317: data = 8'h00;
      17'd45318: data = 8'h00;
      17'd45319: data = 8'h00;
      17'd45320: data = 8'h01;
      17'd45321: data = 8'hfe;
      17'd45322: data = 8'hfe;
      17'd45323: data = 8'h00;
      17'd45324: data = 8'h00;
      17'd45325: data = 8'hfe;
      17'd45326: data = 8'hfe;
      17'd45327: data = 8'hfd;
      17'd45328: data = 8'hfe;
      17'd45329: data = 8'h01;
      17'd45330: data = 8'hfe;
      17'd45331: data = 8'hfe;
      17'd45332: data = 8'hfe;
      17'd45333: data = 8'h00;
      17'd45334: data = 8'h00;
      17'd45335: data = 8'h00;
      17'd45336: data = 8'h00;
      17'd45337: data = 8'h00;
      17'd45338: data = 8'hfd;
      17'd45339: data = 8'hfd;
      17'd45340: data = 8'hfe;
      17'd45341: data = 8'hfe;
      17'd45342: data = 8'hfe;
      17'd45343: data = 8'hfd;
      17'd45344: data = 8'hfc;
      17'd45345: data = 8'h00;
      17'd45346: data = 8'h00;
      17'd45347: data = 8'h00;
      17'd45348: data = 8'h01;
      17'd45349: data = 8'h00;
      17'd45350: data = 8'h01;
      17'd45351: data = 8'h01;
      17'd45352: data = 8'h01;
      17'd45353: data = 8'h00;
      17'd45354: data = 8'hfd;
      17'd45355: data = 8'hfe;
      17'd45356: data = 8'h00;
      17'd45357: data = 8'h00;
      17'd45358: data = 8'hfe;
      17'd45359: data = 8'h01;
      17'd45360: data = 8'h01;
      17'd45361: data = 8'h00;
      17'd45362: data = 8'h02;
      17'd45363: data = 8'h01;
      17'd45364: data = 8'h02;
      17'd45365: data = 8'h01;
      17'd45366: data = 8'hfe;
      17'd45367: data = 8'hfe;
      17'd45368: data = 8'h00;
      17'd45369: data = 8'h00;
      17'd45370: data = 8'hfe;
      17'd45371: data = 8'hfd;
      17'd45372: data = 8'hfc;
      17'd45373: data = 8'hfc;
      17'd45374: data = 8'h00;
      17'd45375: data = 8'h01;
      17'd45376: data = 8'h00;
      17'd45377: data = 8'h00;
      17'd45378: data = 8'h01;
      17'd45379: data = 8'h02;
      17'd45380: data = 8'h01;
      17'd45381: data = 8'hfe;
      17'd45382: data = 8'hfc;
      17'd45383: data = 8'hfa;
      17'd45384: data = 8'hfd;
      17'd45385: data = 8'hfe;
      17'd45386: data = 8'hfd;
      17'd45387: data = 8'hfa;
      17'd45388: data = 8'hfa;
      17'd45389: data = 8'hfe;
      17'd45390: data = 8'hfe;
      17'd45391: data = 8'hfe;
      17'd45392: data = 8'hfd;
      17'd45393: data = 8'hfe;
      17'd45394: data = 8'h02;
      17'd45395: data = 8'h01;
      17'd45396: data = 8'hfe;
      17'd45397: data = 8'hfe;
      17'd45398: data = 8'hfe;
      17'd45399: data = 8'hfe;
      17'd45400: data = 8'hfe;
      17'd45401: data = 8'hfd;
      17'd45402: data = 8'hfc;
      17'd45403: data = 8'hfc;
      17'd45404: data = 8'hfe;
      17'd45405: data = 8'hfe;
      17'd45406: data = 8'hfe;
      17'd45407: data = 8'hfd;
      17'd45408: data = 8'hfe;
      17'd45409: data = 8'h00;
      17'd45410: data = 8'h00;
      17'd45411: data = 8'h00;
      17'd45412: data = 8'hfd;
      17'd45413: data = 8'h00;
      17'd45414: data = 8'hfe;
      17'd45415: data = 8'hfd;
      17'd45416: data = 8'hfe;
      17'd45417: data = 8'hfd;
      17'd45418: data = 8'hfd;
      17'd45419: data = 8'hfd;
      17'd45420: data = 8'hfe;
      17'd45421: data = 8'hfe;
      17'd45422: data = 8'hfe;
      17'd45423: data = 8'h00;
      17'd45424: data = 8'h00;
      17'd45425: data = 8'h01;
      17'd45426: data = 8'h00;
      17'd45427: data = 8'hfe;
      17'd45428: data = 8'h00;
      17'd45429: data = 8'h00;
      17'd45430: data = 8'h00;
      17'd45431: data = 8'h00;
      17'd45432: data = 8'hfd;
      17'd45433: data = 8'hfe;
      17'd45434: data = 8'hfe;
      17'd45435: data = 8'hfe;
      17'd45436: data = 8'h00;
      17'd45437: data = 8'h00;
      17'd45438: data = 8'hfd;
      17'd45439: data = 8'hfe;
      17'd45440: data = 8'h00;
      17'd45441: data = 8'h00;
      17'd45442: data = 8'h00;
      17'd45443: data = 8'h01;
      17'd45444: data = 8'h01;
      17'd45445: data = 8'h00;
      17'd45446: data = 8'h00;
      17'd45447: data = 8'h00;
      17'd45448: data = 8'hfe;
      17'd45449: data = 8'hfe;
      17'd45450: data = 8'hfe;
      17'd45451: data = 8'hfe;
      17'd45452: data = 8'hfd;
      17'd45453: data = 8'hfd;
      17'd45454: data = 8'h00;
      17'd45455: data = 8'hfe;
      17'd45456: data = 8'hfd;
      17'd45457: data = 8'hfe;
      17'd45458: data = 8'h01;
      17'd45459: data = 8'h01;
      17'd45460: data = 8'h00;
      17'd45461: data = 8'h00;
      17'd45462: data = 8'h00;
      17'd45463: data = 8'h00;
      17'd45464: data = 8'h01;
      17'd45465: data = 8'hfe;
      17'd45466: data = 8'hfc;
      17'd45467: data = 8'hfd;
      17'd45468: data = 8'hfe;
      17'd45469: data = 8'h00;
      17'd45470: data = 8'hfe;
      17'd45471: data = 8'hfe;
      17'd45472: data = 8'hfe;
      17'd45473: data = 8'h00;
      17'd45474: data = 8'h01;
      17'd45475: data = 8'h01;
      17'd45476: data = 8'hfe;
      17'd45477: data = 8'hfd;
      17'd45478: data = 8'h00;
      17'd45479: data = 8'h01;
      17'd45480: data = 8'h00;
      17'd45481: data = 8'hfe;
      17'd45482: data = 8'hfe;
      17'd45483: data = 8'h01;
      17'd45484: data = 8'h00;
      17'd45485: data = 8'h00;
      17'd45486: data = 8'hfe;
      17'd45487: data = 8'h00;
      17'd45488: data = 8'h00;
      17'd45489: data = 8'hfe;
      17'd45490: data = 8'h00;
      17'd45491: data = 8'h00;
      17'd45492: data = 8'h00;
      17'd45493: data = 8'h01;
      17'd45494: data = 8'h00;
      17'd45495: data = 8'h00;
      17'd45496: data = 8'h00;
      17'd45497: data = 8'h02;
      17'd45498: data = 8'h04;
      17'd45499: data = 8'h00;
      17'd45500: data = 8'h00;
      17'd45501: data = 8'h01;
      17'd45502: data = 8'h02;
      17'd45503: data = 8'h01;
      17'd45504: data = 8'h00;
      17'd45505: data = 8'h00;
      17'd45506: data = 8'h00;
      17'd45507: data = 8'h02;
      17'd45508: data = 8'h01;
      17'd45509: data = 8'h00;
      17'd45510: data = 8'h00;
      17'd45511: data = 8'h00;
      17'd45512: data = 8'h00;
      17'd45513: data = 8'h01;
      17'd45514: data = 8'hfd;
      17'd45515: data = 8'h00;
      17'd45516: data = 8'h01;
      17'd45517: data = 8'h00;
      17'd45518: data = 8'h01;
      17'd45519: data = 8'h01;
      17'd45520: data = 8'h00;
      17'd45521: data = 8'h00;
      17'd45522: data = 8'h01;
      17'd45523: data = 8'h00;
      17'd45524: data = 8'h01;
      17'd45525: data = 8'h02;
      17'd45526: data = 8'h01;
      17'd45527: data = 8'h00;
      17'd45528: data = 8'hfe;
      17'd45529: data = 8'hfe;
      17'd45530: data = 8'h00;
      17'd45531: data = 8'h00;
      17'd45532: data = 8'h00;
      17'd45533: data = 8'hfe;
      17'd45534: data = 8'h00;
      17'd45535: data = 8'h01;
      17'd45536: data = 8'h01;
      17'd45537: data = 8'h00;
      17'd45538: data = 8'hfe;
      17'd45539: data = 8'h01;
      17'd45540: data = 8'h01;
      17'd45541: data = 8'h01;
      17'd45542: data = 8'h00;
      17'd45543: data = 8'hfe;
      17'd45544: data = 8'hfd;
      17'd45545: data = 8'hfe;
      17'd45546: data = 8'h00;
      17'd45547: data = 8'hfd;
      17'd45548: data = 8'hfd;
      17'd45549: data = 8'hfe;
      17'd45550: data = 8'hfe;
      17'd45551: data = 8'h00;
      17'd45552: data = 8'h00;
      17'd45553: data = 8'hfe;
      17'd45554: data = 8'h00;
      17'd45555: data = 8'h02;
      17'd45556: data = 8'h02;
      17'd45557: data = 8'hfe;
      17'd45558: data = 8'hfe;
      17'd45559: data = 8'hfe;
      17'd45560: data = 8'hfe;
      17'd45561: data = 8'h00;
      17'd45562: data = 8'h00;
      17'd45563: data = 8'hfd;
      17'd45564: data = 8'hfe;
      17'd45565: data = 8'h00;
      17'd45566: data = 8'hfe;
      17'd45567: data = 8'hfe;
      17'd45568: data = 8'hfe;
      17'd45569: data = 8'h00;
      17'd45570: data = 8'h00;
      17'd45571: data = 8'hfe;
      17'd45572: data = 8'hfd;
      17'd45573: data = 8'hfd;
      17'd45574: data = 8'hfe;
      17'd45575: data = 8'hfe;
      17'd45576: data = 8'hfe;
      17'd45577: data = 8'hfd;
      17'd45578: data = 8'hfe;
      17'd45579: data = 8'h00;
      17'd45580: data = 8'h01;
      17'd45581: data = 8'h00;
      17'd45582: data = 8'h00;
      17'd45583: data = 8'hfe;
      17'd45584: data = 8'h00;
      17'd45585: data = 8'h01;
      17'd45586: data = 8'hfe;
      17'd45587: data = 8'hfd;
      17'd45588: data = 8'hfc;
      17'd45589: data = 8'hfd;
      17'd45590: data = 8'hfd;
      17'd45591: data = 8'hfd;
      17'd45592: data = 8'hfd;
      17'd45593: data = 8'hfc;
      17'd45594: data = 8'hfe;
      17'd45595: data = 8'h00;
      17'd45596: data = 8'h01;
      17'd45597: data = 8'hfe;
      17'd45598: data = 8'h00;
      17'd45599: data = 8'h00;
      17'd45600: data = 8'hfe;
      17'd45601: data = 8'hfe;
      17'd45602: data = 8'hfe;
      17'd45603: data = 8'hfd;
      17'd45604: data = 8'hfd;
      17'd45605: data = 8'hfe;
      17'd45606: data = 8'hfe;
      17'd45607: data = 8'hfe;
      17'd45608: data = 8'hfe;
      17'd45609: data = 8'hfd;
      17'd45610: data = 8'hfd;
      17'd45611: data = 8'hfe;
      17'd45612: data = 8'h00;
      17'd45613: data = 8'h00;
      17'd45614: data = 8'hfe;
      17'd45615: data = 8'hfe;
      17'd45616: data = 8'hfd;
      17'd45617: data = 8'hfd;
      17'd45618: data = 8'h00;
      17'd45619: data = 8'hfe;
      17'd45620: data = 8'hfd;
      17'd45621: data = 8'hfe;
      17'd45622: data = 8'hfe;
      17'd45623: data = 8'hfe;
      17'd45624: data = 8'hfe;
      17'd45625: data = 8'h00;
      17'd45626: data = 8'hfe;
      17'd45627: data = 8'hfd;
      17'd45628: data = 8'hfe;
      17'd45629: data = 8'h00;
      17'd45630: data = 8'hfd;
      17'd45631: data = 8'hfe;
      17'd45632: data = 8'hfe;
      17'd45633: data = 8'hfe;
      17'd45634: data = 8'hfd;
      17'd45635: data = 8'hfd;
      17'd45636: data = 8'hfe;
      17'd45637: data = 8'hfe;
      17'd45638: data = 8'hfe;
      17'd45639: data = 8'hfc;
      17'd45640: data = 8'hfd;
      17'd45641: data = 8'hfe;
      17'd45642: data = 8'hfd;
      17'd45643: data = 8'hfe;
      17'd45644: data = 8'hfe;
      17'd45645: data = 8'hfe;
      17'd45646: data = 8'h00;
      17'd45647: data = 8'hfd;
      17'd45648: data = 8'hfe;
      17'd45649: data = 8'hfe;
      17'd45650: data = 8'hfd;
      17'd45651: data = 8'hfd;
      17'd45652: data = 8'hfc;
      17'd45653: data = 8'hfe;
      17'd45654: data = 8'hfd;
      17'd45655: data = 8'hfc;
      17'd45656: data = 8'hfd;
      17'd45657: data = 8'hfd;
      17'd45658: data = 8'hfe;
      17'd45659: data = 8'hfe;
      17'd45660: data = 8'hfe;
      17'd45661: data = 8'h00;
      17'd45662: data = 8'h00;
      17'd45663: data = 8'hfe;
      17'd45664: data = 8'h01;
      17'd45665: data = 8'h00;
      17'd45666: data = 8'h00;
      17'd45667: data = 8'h00;
      17'd45668: data = 8'hfe;
      17'd45669: data = 8'hfe;
      17'd45670: data = 8'hfe;
      17'd45671: data = 8'h00;
      17'd45672: data = 8'hfe;
      17'd45673: data = 8'hfd;
      17'd45674: data = 8'hfe;
      17'd45675: data = 8'h00;
      17'd45676: data = 8'h00;
      17'd45677: data = 8'h00;
      17'd45678: data = 8'hfe;
      17'd45679: data = 8'hfe;
      17'd45680: data = 8'h00;
      17'd45681: data = 8'h00;
      17'd45682: data = 8'hfe;
      17'd45683: data = 8'hfe;
      17'd45684: data = 8'hfe;
      17'd45685: data = 8'hfd;
      17'd45686: data = 8'hfe;
      17'd45687: data = 8'hfd;
      17'd45688: data = 8'hfc;
      17'd45689: data = 8'hfd;
      17'd45690: data = 8'hfd;
      17'd45691: data = 8'hfd;
      17'd45692: data = 8'hfd;
      17'd45693: data = 8'hfd;
      17'd45694: data = 8'hfc;
      17'd45695: data = 8'hfc;
      17'd45696: data = 8'hfa;
      17'd45697: data = 8'hfd;
      17'd45698: data = 8'hfc;
      17'd45699: data = 8'hfd;
      17'd45700: data = 8'hfd;
      17'd45701: data = 8'hfd;
      17'd45702: data = 8'hfe;
      17'd45703: data = 8'hfd;
      17'd45704: data = 8'hfe;
      17'd45705: data = 8'hfd;
      17'd45706: data = 8'hfe;
      17'd45707: data = 8'h01;
      17'd45708: data = 8'hfe;
      17'd45709: data = 8'hfe;
      17'd45710: data = 8'hfe;
      17'd45711: data = 8'hfe;
      17'd45712: data = 8'hfe;
      17'd45713: data = 8'hfe;
      17'd45714: data = 8'hfe;
      17'd45715: data = 8'hfe;
      17'd45716: data = 8'hfd;
      17'd45717: data = 8'hfc;
      17'd45718: data = 8'hfd;
      17'd45719: data = 8'h00;
      17'd45720: data = 8'hfe;
      17'd45721: data = 8'hfe;
      17'd45722: data = 8'hfe;
      17'd45723: data = 8'hfe;
      17'd45724: data = 8'h00;
      17'd45725: data = 8'h00;
      17'd45726: data = 8'hfe;
      17'd45727: data = 8'hfe;
      17'd45728: data = 8'hfe;
      17'd45729: data = 8'h00;
      17'd45730: data = 8'h00;
      17'd45731: data = 8'hfe;
      17'd45732: data = 8'h00;
      17'd45733: data = 8'hfe;
      17'd45734: data = 8'hfe;
      17'd45735: data = 8'h00;
      17'd45736: data = 8'h00;
      17'd45737: data = 8'h00;
      17'd45738: data = 8'h01;
      17'd45739: data = 8'h02;
      17'd45740: data = 8'h00;
      17'd45741: data = 8'h00;
      17'd45742: data = 8'hfe;
      17'd45743: data = 8'hfe;
      17'd45744: data = 8'h00;
      17'd45745: data = 8'hfe;
      17'd45746: data = 8'hfd;
      17'd45747: data = 8'hfd;
      17'd45748: data = 8'hfd;
      17'd45749: data = 8'hfe;
      17'd45750: data = 8'h00;
      17'd45751: data = 8'hfe;
      17'd45752: data = 8'hfe;
      17'd45753: data = 8'h00;
      17'd45754: data = 8'h02;
      17'd45755: data = 8'h04;
      17'd45756: data = 8'h01;
      17'd45757: data = 8'h00;
      17'd45758: data = 8'h01;
      17'd45759: data = 8'h02;
      17'd45760: data = 8'h02;
      17'd45761: data = 8'h00;
      17'd45762: data = 8'h00;
      17'd45763: data = 8'h00;
      17'd45764: data = 8'h00;
      17'd45765: data = 8'h00;
      17'd45766: data = 8'hfe;
      17'd45767: data = 8'h00;
      17'd45768: data = 8'h01;
      17'd45769: data = 8'h00;
      17'd45770: data = 8'h00;
      17'd45771: data = 8'h01;
      17'd45772: data = 8'h01;
      17'd45773: data = 8'h02;
      17'd45774: data = 8'h02;
      17'd45775: data = 8'h00;
      17'd45776: data = 8'hfe;
      17'd45777: data = 8'h01;
      17'd45778: data = 8'h00;
      17'd45779: data = 8'hfe;
      17'd45780: data = 8'hfe;
      17'd45781: data = 8'hfe;
      17'd45782: data = 8'h00;
      17'd45783: data = 8'h00;
      17'd45784: data = 8'h00;
      17'd45785: data = 8'hfd;
      17'd45786: data = 8'hfd;
      17'd45787: data = 8'h00;
      17'd45788: data = 8'hfe;
      17'd45789: data = 8'hfe;
      17'd45790: data = 8'hfe;
      17'd45791: data = 8'h00;
      17'd45792: data = 8'h00;
      17'd45793: data = 8'h00;
      17'd45794: data = 8'h01;
      17'd45795: data = 8'h01;
      17'd45796: data = 8'hfd;
      17'd45797: data = 8'h00;
      17'd45798: data = 8'h00;
      17'd45799: data = 8'h00;
      17'd45800: data = 8'h00;
      17'd45801: data = 8'h00;
      17'd45802: data = 8'h00;
      17'd45803: data = 8'h00;
      17'd45804: data = 8'h00;
      17'd45805: data = 8'h00;
      17'd45806: data = 8'h00;
      17'd45807: data = 8'h01;
      17'd45808: data = 8'h01;
      17'd45809: data = 8'h01;
      17'd45810: data = 8'h00;
      17'd45811: data = 8'h01;
      17'd45812: data = 8'h00;
      17'd45813: data = 8'h00;
      17'd45814: data = 8'h00;
      17'd45815: data = 8'h01;
      17'd45816: data = 8'hfe;
      17'd45817: data = 8'hfd;
      17'd45818: data = 8'hfd;
      17'd45819: data = 8'hfd;
      17'd45820: data = 8'hfe;
      17'd45821: data = 8'hfe;
      17'd45822: data = 8'hfe;
      17'd45823: data = 8'h00;
      17'd45824: data = 8'hfe;
      17'd45825: data = 8'h00;
      17'd45826: data = 8'h00;
      17'd45827: data = 8'h00;
      17'd45828: data = 8'h01;
      17'd45829: data = 8'h01;
      17'd45830: data = 8'hfe;
      17'd45831: data = 8'hfe;
      17'd45832: data = 8'hfd;
      17'd45833: data = 8'hfc;
      17'd45834: data = 8'hfd;
      17'd45835: data = 8'hfe;
      17'd45836: data = 8'hfe;
      17'd45837: data = 8'hfd;
      17'd45838: data = 8'hfc;
      17'd45839: data = 8'hfc;
      17'd45840: data = 8'hfe;
      17'd45841: data = 8'h00;
      17'd45842: data = 8'hfe;
      17'd45843: data = 8'hfe;
      17'd45844: data = 8'h00;
      17'd45845: data = 8'hfe;
      17'd45846: data = 8'h00;
      17'd45847: data = 8'hfe;
      17'd45848: data = 8'hfe;
      17'd45849: data = 8'hfd;
      17'd45850: data = 8'hfe;
      17'd45851: data = 8'h01;
      17'd45852: data = 8'hfe;
      17'd45853: data = 8'h01;
      17'd45854: data = 8'h00;
      17'd45855: data = 8'hfe;
      17'd45856: data = 8'h01;
      17'd45857: data = 8'h02;
      17'd45858: data = 8'h00;
      17'd45859: data = 8'hfe;
      17'd45860: data = 8'h00;
      17'd45861: data = 8'h00;
      17'd45862: data = 8'h01;
      17'd45863: data = 8'h00;
      17'd45864: data = 8'h00;
      17'd45865: data = 8'hfe;
      17'd45866: data = 8'hfe;
      17'd45867: data = 8'h01;
      17'd45868: data = 8'h01;
      17'd45869: data = 8'h00;
      17'd45870: data = 8'h01;
      17'd45871: data = 8'h00;
      17'd45872: data = 8'h00;
      17'd45873: data = 8'h00;
      17'd45874: data = 8'h01;
      17'd45875: data = 8'h00;
      17'd45876: data = 8'hfe;
      17'd45877: data = 8'hfe;
      17'd45878: data = 8'hfe;
      17'd45879: data = 8'hfd;
      17'd45880: data = 8'h00;
      17'd45881: data = 8'h01;
      17'd45882: data = 8'hfe;
      17'd45883: data = 8'hfe;
      17'd45884: data = 8'h00;
      17'd45885: data = 8'h01;
      17'd45886: data = 8'h01;
      17'd45887: data = 8'h00;
      17'd45888: data = 8'hfe;
      17'd45889: data = 8'h00;
      17'd45890: data = 8'hfe;
      17'd45891: data = 8'h00;
      17'd45892: data = 8'hfe;
      17'd45893: data = 8'hfd;
      17'd45894: data = 8'hfd;
      17'd45895: data = 8'hfd;
      17'd45896: data = 8'hfe;
      17'd45897: data = 8'hfe;
      17'd45898: data = 8'hfe;
      17'd45899: data = 8'hfe;
      17'd45900: data = 8'hfe;
      17'd45901: data = 8'h00;
      17'd45902: data = 8'h02;
      17'd45903: data = 8'h01;
      17'd45904: data = 8'h00;
      17'd45905: data = 8'h01;
      17'd45906: data = 8'h00;
      17'd45907: data = 8'h00;
      17'd45908: data = 8'hfe;
      17'd45909: data = 8'hfe;
      17'd45910: data = 8'hfe;
      17'd45911: data = 8'h00;
      17'd45912: data = 8'h01;
      17'd45913: data = 8'h00;
      17'd45914: data = 8'h00;
      17'd45915: data = 8'hfe;
      17'd45916: data = 8'h00;
      17'd45917: data = 8'h01;
      17'd45918: data = 8'h00;
      17'd45919: data = 8'hfe;
      17'd45920: data = 8'hfe;
      17'd45921: data = 8'h00;
      17'd45922: data = 8'h01;
      17'd45923: data = 8'h00;
      17'd45924: data = 8'h00;
      17'd45925: data = 8'hfe;
      17'd45926: data = 8'h00;
      17'd45927: data = 8'h02;
      17'd45928: data = 8'h00;
      17'd45929: data = 8'h00;
      17'd45930: data = 8'h01;
      17'd45931: data = 8'h01;
      17'd45932: data = 8'h01;
      17'd45933: data = 8'h02;
      17'd45934: data = 8'h01;
      17'd45935: data = 8'h02;
      17'd45936: data = 8'h00;
      17'd45937: data = 8'hfe;
      17'd45938: data = 8'h01;
      17'd45939: data = 8'h00;
      17'd45940: data = 8'h00;
      17'd45941: data = 8'h00;
      17'd45942: data = 8'h00;
      17'd45943: data = 8'hfe;
      17'd45944: data = 8'hfe;
      17'd45945: data = 8'h01;
      17'd45946: data = 8'h00;
      17'd45947: data = 8'hfd;
      17'd45948: data = 8'hfd;
      17'd45949: data = 8'hfe;
      17'd45950: data = 8'h00;
      17'd45951: data = 8'hfe;
      17'd45952: data = 8'hfd;
      17'd45953: data = 8'hfd;
      17'd45954: data = 8'hfe;
      17'd45955: data = 8'h00;
      17'd45956: data = 8'hfe;
      17'd45957: data = 8'hfd;
      17'd45958: data = 8'hfc;
      17'd45959: data = 8'hfe;
      17'd45960: data = 8'h00;
      17'd45961: data = 8'hfd;
      17'd45962: data = 8'hfd;
      17'd45963: data = 8'hfc;
      17'd45964: data = 8'hfd;
      17'd45965: data = 8'hfe;
      17'd45966: data = 8'h00;
      17'd45967: data = 8'h00;
      17'd45968: data = 8'hfe;
      17'd45969: data = 8'h00;
      17'd45970: data = 8'h00;
      17'd45971: data = 8'h00;
      17'd45972: data = 8'h00;
      17'd45973: data = 8'hfe;
      17'd45974: data = 8'hfe;
      17'd45975: data = 8'hfe;
      17'd45976: data = 8'hfe;
      17'd45977: data = 8'hfd;
      17'd45978: data = 8'hfd;
      17'd45979: data = 8'hfe;
      17'd45980: data = 8'h00;
      17'd45981: data = 8'h00;
      17'd45982: data = 8'hfe;
      17'd45983: data = 8'hfe;
      17'd45984: data = 8'h00;
      17'd45985: data = 8'h00;
      17'd45986: data = 8'hfe;
      17'd45987: data = 8'hfd;
      17'd45988: data = 8'hfd;
      17'd45989: data = 8'hfe;
      17'd45990: data = 8'hfd;
      17'd45991: data = 8'hfe;
      17'd45992: data = 8'hfd;
      17'd45993: data = 8'hfd;
      17'd45994: data = 8'h00;
      17'd45995: data = 8'h00;
      17'd45996: data = 8'h00;
      17'd45997: data = 8'hfe;
      17'd45998: data = 8'hfe;
      17'd45999: data = 8'h01;
      17'd46000: data = 8'h00;
      17'd46001: data = 8'hfe;
      17'd46002: data = 8'hfe;
      17'd46003: data = 8'hfd;
      17'd46004: data = 8'hfd;
      17'd46005: data = 8'hfe;
      17'd46006: data = 8'hfe;
      17'd46007: data = 8'hfd;
      17'd46008: data = 8'hfc;
      17'd46009: data = 8'hfe;
      17'd46010: data = 8'h00;
      17'd46011: data = 8'h00;
      17'd46012: data = 8'h00;
      17'd46013: data = 8'h00;
      17'd46014: data = 8'h01;
      17'd46015: data = 8'h02;
      17'd46016: data = 8'h01;
      17'd46017: data = 8'hfe;
      17'd46018: data = 8'hfe;
      17'd46019: data = 8'hfe;
      17'd46020: data = 8'hfe;
      17'd46021: data = 8'hfd;
      17'd46022: data = 8'hfe;
      17'd46023: data = 8'hfe;
      17'd46024: data = 8'hfe;
      17'd46025: data = 8'h01;
      17'd46026: data = 8'h01;
      17'd46027: data = 8'h00;
      17'd46028: data = 8'h01;
      17'd46029: data = 8'h01;
      17'd46030: data = 8'h00;
      17'd46031: data = 8'h01;
      17'd46032: data = 8'h01;
      17'd46033: data = 8'h00;
      17'd46034: data = 8'hfe;
      17'd46035: data = 8'h00;
      17'd46036: data = 8'h00;
      17'd46037: data = 8'hfd;
      17'd46038: data = 8'hfd;
      17'd46039: data = 8'hfe;
      17'd46040: data = 8'h00;
      17'd46041: data = 8'h01;
      17'd46042: data = 8'h01;
      17'd46043: data = 8'h01;
      17'd46044: data = 8'h01;
      17'd46045: data = 8'h01;
      17'd46046: data = 8'h00;
      17'd46047: data = 8'h00;
      17'd46048: data = 8'hfe;
      17'd46049: data = 8'hfd;
      17'd46050: data = 8'hfd;
      17'd46051: data = 8'hfe;
      17'd46052: data = 8'hfe;
      17'd46053: data = 8'h00;
      17'd46054: data = 8'h01;
      17'd46055: data = 8'h00;
      17'd46056: data = 8'h00;
      17'd46057: data = 8'h00;
      17'd46058: data = 8'h00;
      17'd46059: data = 8'hfe;
      17'd46060: data = 8'hfe;
      17'd46061: data = 8'h00;
      17'd46062: data = 8'h00;
      17'd46063: data = 8'h00;
      17'd46064: data = 8'hfe;
      17'd46065: data = 8'h00;
      17'd46066: data = 8'h00;
      17'd46067: data = 8'hfe;
      17'd46068: data = 8'h00;
      17'd46069: data = 8'h00;
      17'd46070: data = 8'h00;
      17'd46071: data = 8'h00;
      17'd46072: data = 8'h01;
      17'd46073: data = 8'h01;
      17'd46074: data = 8'h00;
      17'd46075: data = 8'h00;
      17'd46076: data = 8'hfe;
      17'd46077: data = 8'hfd;
      17'd46078: data = 8'hfd;
      17'd46079: data = 8'hfd;
      17'd46080: data = 8'hfd;
      17'd46081: data = 8'hfd;
      17'd46082: data = 8'hfe;
      17'd46083: data = 8'hfe;
      17'd46084: data = 8'h00;
      17'd46085: data = 8'h00;
      17'd46086: data = 8'h00;
      17'd46087: data = 8'h01;
      17'd46088: data = 8'h01;
      17'd46089: data = 8'hfe;
      17'd46090: data = 8'hfe;
      17'd46091: data = 8'hfe;
      17'd46092: data = 8'hfd;
      17'd46093: data = 8'hfe;
      17'd46094: data = 8'hfe;
      17'd46095: data = 8'hfe;
      17'd46096: data = 8'h00;
      17'd46097: data = 8'h00;
      17'd46098: data = 8'hfe;
      17'd46099: data = 8'h01;
      17'd46100: data = 8'h00;
      17'd46101: data = 8'h00;
      17'd46102: data = 8'h02;
      17'd46103: data = 8'h02;
      17'd46104: data = 8'h01;
      17'd46105: data = 8'h00;
      17'd46106: data = 8'h00;
      17'd46107: data = 8'h00;
      17'd46108: data = 8'h00;
      17'd46109: data = 8'h00;
      17'd46110: data = 8'h00;
      17'd46111: data = 8'h00;
      17'd46112: data = 8'h00;
      17'd46113: data = 8'h01;
      17'd46114: data = 8'h00;
      17'd46115: data = 8'h01;
      17'd46116: data = 8'h01;
      17'd46117: data = 8'h01;
      17'd46118: data = 8'h00;
      17'd46119: data = 8'h00;
      17'd46120: data = 8'h00;
      17'd46121: data = 8'hfe;
      17'd46122: data = 8'h00;
      17'd46123: data = 8'hfe;
      17'd46124: data = 8'h00;
      17'd46125: data = 8'h00;
      17'd46126: data = 8'h00;
      17'd46127: data = 8'h01;
      17'd46128: data = 8'h00;
      17'd46129: data = 8'h00;
      17'd46130: data = 8'h01;
      17'd46131: data = 8'h00;
      17'd46132: data = 8'h00;
      17'd46133: data = 8'h01;
      17'd46134: data = 8'hfe;
      17'd46135: data = 8'hfe;
      17'd46136: data = 8'hfd;
      17'd46137: data = 8'hfd;
      17'd46138: data = 8'hfe;
      17'd46139: data = 8'hfe;
      17'd46140: data = 8'hfe;
      17'd46141: data = 8'hfe;
      17'd46142: data = 8'h01;
      17'd46143: data = 8'h01;
      17'd46144: data = 8'h00;
      17'd46145: data = 8'h00;
      17'd46146: data = 8'h01;
      17'd46147: data = 8'h00;
      17'd46148: data = 8'hfe;
      17'd46149: data = 8'hfe;
      17'd46150: data = 8'hfe;
      17'd46151: data = 8'hfd;
      17'd46152: data = 8'hfe;
      17'd46153: data = 8'hfd;
      17'd46154: data = 8'h00;
      17'd46155: data = 8'h01;
      17'd46156: data = 8'h00;
      17'd46157: data = 8'h01;
      17'd46158: data = 8'h02;
      17'd46159: data = 8'h01;
      17'd46160: data = 8'h01;
      17'd46161: data = 8'h00;
      17'd46162: data = 8'h01;
      17'd46163: data = 8'h01;
      17'd46164: data = 8'hfe;
      17'd46165: data = 8'hfd;
      17'd46166: data = 8'hfd;
      17'd46167: data = 8'hfe;
      17'd46168: data = 8'hfe;
      17'd46169: data = 8'hfe;
      17'd46170: data = 8'hfe;
      17'd46171: data = 8'h00;
      17'd46172: data = 8'h00;
      17'd46173: data = 8'h01;
      17'd46174: data = 8'hfe;
      17'd46175: data = 8'h00;
      17'd46176: data = 8'h01;
      17'd46177: data = 8'hfe;
      17'd46178: data = 8'hfe;
      17'd46179: data = 8'hfe;
      17'd46180: data = 8'hfe;
      17'd46181: data = 8'hfe;
      17'd46182: data = 8'hfe;
      17'd46183: data = 8'hfe;
      17'd46184: data = 8'h00;
      17'd46185: data = 8'h00;
      17'd46186: data = 8'hfe;
      17'd46187: data = 8'h01;
      17'd46188: data = 8'h01;
      17'd46189: data = 8'hfe;
      17'd46190: data = 8'hfe;
      17'd46191: data = 8'hfe;
      17'd46192: data = 8'h00;
      17'd46193: data = 8'h00;
      17'd46194: data = 8'hfe;
      17'd46195: data = 8'hfe;
      17'd46196: data = 8'hfe;
      17'd46197: data = 8'h00;
      17'd46198: data = 8'h02;
      17'd46199: data = 8'h00;
      17'd46200: data = 8'h00;
      17'd46201: data = 8'h00;
      17'd46202: data = 8'h01;
      17'd46203: data = 8'h01;
      17'd46204: data = 8'hfe;
      17'd46205: data = 8'hfe;
      17'd46206: data = 8'h00;
      17'd46207: data = 8'h00;
      17'd46208: data = 8'h00;
      17'd46209: data = 8'h00;
      17'd46210: data = 8'hfe;
      17'd46211: data = 8'h00;
      17'd46212: data = 8'hfe;
      17'd46213: data = 8'hfe;
      17'd46214: data = 8'h00;
      17'd46215: data = 8'h00;
      17'd46216: data = 8'hfe;
      17'd46217: data = 8'h00;
      17'd46218: data = 8'h00;
      17'd46219: data = 8'hfe;
      17'd46220: data = 8'hfe;
      17'd46221: data = 8'h00;
      17'd46222: data = 8'h00;
      17'd46223: data = 8'h00;
      17'd46224: data = 8'h01;
      17'd46225: data = 8'h02;
      17'd46226: data = 8'h01;
      17'd46227: data = 8'h01;
      17'd46228: data = 8'h01;
      17'd46229: data = 8'h00;
      17'd46230: data = 8'hfe;
      17'd46231: data = 8'hfe;
      17'd46232: data = 8'hfe;
      17'd46233: data = 8'hfe;
      17'd46234: data = 8'h00;
      17'd46235: data = 8'h01;
      17'd46236: data = 8'h01;
      17'd46237: data = 8'h00;
      17'd46238: data = 8'h01;
      17'd46239: data = 8'h01;
      17'd46240: data = 8'h01;
      17'd46241: data = 8'h01;
      17'd46242: data = 8'h01;
      17'd46243: data = 8'h01;
      17'd46244: data = 8'h01;
      17'd46245: data = 8'h01;
      17'd46246: data = 8'h00;
      17'd46247: data = 8'hfe;
      17'd46248: data = 8'hfd;
      17'd46249: data = 8'hfe;
      17'd46250: data = 8'hfe;
      17'd46251: data = 8'hfd;
      17'd46252: data = 8'hfe;
      17'd46253: data = 8'h00;
      17'd46254: data = 8'h00;
      17'd46255: data = 8'h01;
      17'd46256: data = 8'h01;
      17'd46257: data = 8'h02;
      17'd46258: data = 8'h00;
      17'd46259: data = 8'hfe;
      17'd46260: data = 8'h00;
      17'd46261: data = 8'hfe;
      17'd46262: data = 8'hfd;
      17'd46263: data = 8'hfc;
      17'd46264: data = 8'hfc;
      17'd46265: data = 8'hfd;
      17'd46266: data = 8'hfe;
      17'd46267: data = 8'hfe;
      17'd46268: data = 8'hfe;
      17'd46269: data = 8'hfe;
      17'd46270: data = 8'h00;
      17'd46271: data = 8'h01;
      17'd46272: data = 8'h00;
      17'd46273: data = 8'hfe;
      17'd46274: data = 8'h00;
      17'd46275: data = 8'h01;
      17'd46276: data = 8'h00;
      17'd46277: data = 8'hfe;
      17'd46278: data = 8'hfe;
      17'd46279: data = 8'hfd;
      17'd46280: data = 8'hfd;
      17'd46281: data = 8'hfe;
      17'd46282: data = 8'hfe;
      17'd46283: data = 8'hfe;
      17'd46284: data = 8'h00;
      17'd46285: data = 8'h01;
      17'd46286: data = 8'h01;
      17'd46287: data = 8'h01;
      17'd46288: data = 8'h01;
      17'd46289: data = 8'h00;
      17'd46290: data = 8'h00;
      17'd46291: data = 8'h00;
      17'd46292: data = 8'hfd;
      17'd46293: data = 8'hfe;
      17'd46294: data = 8'hfe;
      17'd46295: data = 8'hfe;
      17'd46296: data = 8'h01;
      17'd46297: data = 8'h00;
      17'd46298: data = 8'h00;
      17'd46299: data = 8'h04;
      17'd46300: data = 8'h02;
      17'd46301: data = 8'h00;
      17'd46302: data = 8'h00;
      17'd46303: data = 8'h02;
      17'd46304: data = 8'h00;
      17'd46305: data = 8'h00;
      17'd46306: data = 8'h00;
      17'd46307: data = 8'hfd;
      17'd46308: data = 8'hfd;
      17'd46309: data = 8'hfe;
      17'd46310: data = 8'h00;
      17'd46311: data = 8'h00;
      17'd46312: data = 8'h01;
      17'd46313: data = 8'h00;
      17'd46314: data = 8'h01;
      17'd46315: data = 8'h04;
      17'd46316: data = 8'h02;
      17'd46317: data = 8'h04;
      17'd46318: data = 8'h02;
      17'd46319: data = 8'h01;
      17'd46320: data = 8'h02;
      17'd46321: data = 8'h00;
      17'd46322: data = 8'h00;
      17'd46323: data = 8'h00;
      17'd46324: data = 8'h00;
      17'd46325: data = 8'h00;
      17'd46326: data = 8'h01;
      17'd46327: data = 8'h00;
      17'd46328: data = 8'h01;
      17'd46329: data = 8'h01;
      17'd46330: data = 8'h01;
      17'd46331: data = 8'h01;
      17'd46332: data = 8'h02;
      17'd46333: data = 8'h02;
      17'd46334: data = 8'h00;
      17'd46335: data = 8'h00;
      17'd46336: data = 8'h01;
      17'd46337: data = 8'h01;
      17'd46338: data = 8'h00;
      17'd46339: data = 8'hfe;
      17'd46340: data = 8'hfe;
      17'd46341: data = 8'h00;
      17'd46342: data = 8'h00;
      17'd46343: data = 8'h00;
      17'd46344: data = 8'h01;
      17'd46345: data = 8'h01;
      17'd46346: data = 8'h00;
      17'd46347: data = 8'h01;
      17'd46348: data = 8'h02;
      17'd46349: data = 8'h00;
      17'd46350: data = 8'hfe;
      17'd46351: data = 8'hfe;
      17'd46352: data = 8'hfe;
      17'd46353: data = 8'h00;
      17'd46354: data = 8'h00;
      17'd46355: data = 8'hfe;
      17'd46356: data = 8'hfe;
      17'd46357: data = 8'h00;
      17'd46358: data = 8'hfe;
      17'd46359: data = 8'h00;
      17'd46360: data = 8'h00;
      17'd46361: data = 8'h00;
      17'd46362: data = 8'h01;
      17'd46363: data = 8'hfe;
      17'd46364: data = 8'h00;
      17'd46365: data = 8'h00;
      17'd46366: data = 8'h00;
      17'd46367: data = 8'h00;
      17'd46368: data = 8'h00;
      17'd46369: data = 8'h00;
      17'd46370: data = 8'h01;
      17'd46371: data = 8'h00;
      17'd46372: data = 8'h00;
      17'd46373: data = 8'h01;
      17'd46374: data = 8'h00;
      17'd46375: data = 8'h00;
      17'd46376: data = 8'h00;
      17'd46377: data = 8'hfe;
      17'd46378: data = 8'hfe;
      17'd46379: data = 8'h00;
      17'd46380: data = 8'hfe;
      17'd46381: data = 8'hfd;
      17'd46382: data = 8'hfd;
      17'd46383: data = 8'h00;
      17'd46384: data = 8'h00;
      17'd46385: data = 8'h00;
      17'd46386: data = 8'h01;
      17'd46387: data = 8'h00;
      17'd46388: data = 8'h00;
      17'd46389: data = 8'h01;
      17'd46390: data = 8'h02;
      17'd46391: data = 8'h00;
      17'd46392: data = 8'hfd;
      17'd46393: data = 8'h00;
      17'd46394: data = 8'h00;
      17'd46395: data = 8'hfe;
      17'd46396: data = 8'hfe;
      17'd46397: data = 8'hfe;
      17'd46398: data = 8'hfd;
      17'd46399: data = 8'hfe;
      17'd46400: data = 8'h01;
      17'd46401: data = 8'hfe;
      17'd46402: data = 8'h00;
      17'd46403: data = 8'h01;
      17'd46404: data = 8'h00;
      17'd46405: data = 8'h00;
      17'd46406: data = 8'hfe;
      17'd46407: data = 8'hfe;
      17'd46408: data = 8'hfe;
      17'd46409: data = 8'hfe;
      17'd46410: data = 8'h00;
      17'd46411: data = 8'hfe;
      17'd46412: data = 8'hfe;
      17'd46413: data = 8'hfe;
      17'd46414: data = 8'h00;
      17'd46415: data = 8'hfe;
      17'd46416: data = 8'h00;
      17'd46417: data = 8'h01;
      17'd46418: data = 8'h01;
      17'd46419: data = 8'h01;
      17'd46420: data = 8'h02;
      17'd46421: data = 8'h01;
      17'd46422: data = 8'h00;
      17'd46423: data = 8'h01;
      17'd46424: data = 8'hfe;
      17'd46425: data = 8'hfd;
      17'd46426: data = 8'hfe;
      17'd46427: data = 8'hfe;
      17'd46428: data = 8'hfe;
      17'd46429: data = 8'hfe;
      17'd46430: data = 8'hfe;
      17'd46431: data = 8'h00;
      17'd46432: data = 8'h01;
      17'd46433: data = 8'h00;
      17'd46434: data = 8'h00;
      17'd46435: data = 8'hfe;
      17'd46436: data = 8'hfe;
      17'd46437: data = 8'hfe;
      17'd46438: data = 8'hfe;
      17'd46439: data = 8'hfe;
      17'd46440: data = 8'hfc;
      17'd46441: data = 8'hfc;
      17'd46442: data = 8'hfd;
      17'd46443: data = 8'hfe;
      17'd46444: data = 8'hfe;
      17'd46445: data = 8'hfe;
      17'd46446: data = 8'hfe;
      17'd46447: data = 8'h00;
      17'd46448: data = 8'h00;
      17'd46449: data = 8'hfe;
      17'd46450: data = 8'h00;
      17'd46451: data = 8'h00;
      17'd46452: data = 8'hfe;
      17'd46453: data = 8'hfe;
      17'd46454: data = 8'hfe;
      17'd46455: data = 8'hfe;
      17'd46456: data = 8'hfe;
      17'd46457: data = 8'hfe;
      17'd46458: data = 8'hfe;
      17'd46459: data = 8'hfe;
      17'd46460: data = 8'hfe;
      17'd46461: data = 8'hfd;
      17'd46462: data = 8'hfe;
      17'd46463: data = 8'h00;
      17'd46464: data = 8'h00;
      17'd46465: data = 8'h00;
      17'd46466: data = 8'hfe;
      17'd46467: data = 8'h00;
      17'd46468: data = 8'hfe;
      17'd46469: data = 8'hfe;
      17'd46470: data = 8'hfc;
      17'd46471: data = 8'hfc;
      17'd46472: data = 8'hfe;
      17'd46473: data = 8'hfc;
      17'd46474: data = 8'hfc;
      17'd46475: data = 8'hfd;
      17'd46476: data = 8'hfd;
      17'd46477: data = 8'hfd;
      17'd46478: data = 8'hfe;
      17'd46479: data = 8'h00;
      17'd46480: data = 8'hfe;
      17'd46481: data = 8'h00;
      17'd46482: data = 8'h00;
      17'd46483: data = 8'hfe;
      17'd46484: data = 8'hfd;
      17'd46485: data = 8'hfe;
      17'd46486: data = 8'hfe;
      17'd46487: data = 8'hfe;
      17'd46488: data = 8'h00;
      17'd46489: data = 8'h00;
      17'd46490: data = 8'h00;
      17'd46491: data = 8'h00;
      17'd46492: data = 8'hfe;
      17'd46493: data = 8'h00;
      17'd46494: data = 8'h01;
      17'd46495: data = 8'h01;
      17'd46496: data = 8'h00;
      17'd46497: data = 8'h00;
      17'd46498: data = 8'h01;
      17'd46499: data = 8'hfe;
      17'd46500: data = 8'hfe;
      17'd46501: data = 8'hfe;
      17'd46502: data = 8'hfe;
      17'd46503: data = 8'hfe;
      17'd46504: data = 8'hfe;
      17'd46505: data = 8'hfe;
      17'd46506: data = 8'hfe;
      17'd46507: data = 8'hfe;
      17'd46508: data = 8'hfe;
      17'd46509: data = 8'h00;
      17'd46510: data = 8'h00;
      17'd46511: data = 8'h02;
      17'd46512: data = 8'hfe;
      17'd46513: data = 8'hfd;
      17'd46514: data = 8'hfe;
      17'd46515: data = 8'hfe;
      17'd46516: data = 8'h00;
      17'd46517: data = 8'h00;
      17'd46518: data = 8'hfe;
      17'd46519: data = 8'hfe;
      17'd46520: data = 8'h00;
      17'd46521: data = 8'h00;
      17'd46522: data = 8'h01;
      17'd46523: data = 8'hfd;
      17'd46524: data = 8'hfe;
      17'd46525: data = 8'hfe;
      17'd46526: data = 8'hfe;
      17'd46527: data = 8'hfe;
      17'd46528: data = 8'hfe;
      17'd46529: data = 8'hfe;
      17'd46530: data = 8'h00;
      17'd46531: data = 8'hfe;
      17'd46532: data = 8'hfe;
      17'd46533: data = 8'hfd;
      17'd46534: data = 8'hfe;
      17'd46535: data = 8'hfe;
      17'd46536: data = 8'hfe;
      17'd46537: data = 8'hfe;
      17'd46538: data = 8'h00;
      17'd46539: data = 8'h00;
      17'd46540: data = 8'h00;
      17'd46541: data = 8'h00;
      17'd46542: data = 8'hfe;
      17'd46543: data = 8'h00;
      17'd46544: data = 8'h00;
      17'd46545: data = 8'h00;
      17'd46546: data = 8'h00;
      17'd46547: data = 8'hfe;
      17'd46548: data = 8'hfe;
      17'd46549: data = 8'h00;
      17'd46550: data = 8'hfe;
      17'd46551: data = 8'h00;
      17'd46552: data = 8'hfe;
      17'd46553: data = 8'hfe;
      17'd46554: data = 8'h00;
      17'd46555: data = 8'h00;
      17'd46556: data = 8'h01;
      17'd46557: data = 8'hfe;
      17'd46558: data = 8'h00;
      17'd46559: data = 8'h00;
      17'd46560: data = 8'hfe;
      17'd46561: data = 8'hfe;
      17'd46562: data = 8'hfe;
      17'd46563: data = 8'h00;
      17'd46564: data = 8'hfe;
      17'd46565: data = 8'hfe;
      17'd46566: data = 8'hfe;
      17'd46567: data = 8'hfe;
      17'd46568: data = 8'hfe;
      17'd46569: data = 8'h00;
      17'd46570: data = 8'hfe;
      17'd46571: data = 8'hfe;
      17'd46572: data = 8'h01;
      17'd46573: data = 8'h00;
      17'd46574: data = 8'hfd;
      17'd46575: data = 8'hfd;
      17'd46576: data = 8'hfe;
      17'd46577: data = 8'hfe;
      17'd46578: data = 8'hfd;
      17'd46579: data = 8'hfd;
      17'd46580: data = 8'hfc;
      17'd46581: data = 8'hfd;
      17'd46582: data = 8'hfd;
      17'd46583: data = 8'hfe;
      17'd46584: data = 8'hfe;
      17'd46585: data = 8'hfe;
      17'd46586: data = 8'hfd;
      17'd46587: data = 8'hfe;
      17'd46588: data = 8'h00;
      17'd46589: data = 8'h00;
      17'd46590: data = 8'hfe;
      17'd46591: data = 8'hfe;
      17'd46592: data = 8'h00;
      17'd46593: data = 8'hfe;
      17'd46594: data = 8'hfe;
      17'd46595: data = 8'hfe;
      17'd46596: data = 8'hfd;
      17'd46597: data = 8'hfd;
      17'd46598: data = 8'hfd;
      17'd46599: data = 8'hfe;
      17'd46600: data = 8'h00;
      17'd46601: data = 8'h00;
      17'd46602: data = 8'h00;
      17'd46603: data = 8'h00;
      17'd46604: data = 8'h00;
      17'd46605: data = 8'h00;
      17'd46606: data = 8'hfe;
      17'd46607: data = 8'h00;
      17'd46608: data = 8'hfe;
      17'd46609: data = 8'hfd;
      17'd46610: data = 8'hfd;
      17'd46611: data = 8'hfd;
      17'd46612: data = 8'hfe;
      17'd46613: data = 8'hfd;
      17'd46614: data = 8'hfe;
      17'd46615: data = 8'hfd;
      17'd46616: data = 8'h00;
      17'd46617: data = 8'h00;
      17'd46618: data = 8'h00;
      17'd46619: data = 8'hfe;
      17'd46620: data = 8'h00;
      17'd46621: data = 8'h02;
      17'd46622: data = 8'hfe;
      17'd46623: data = 8'h00;
      17'd46624: data = 8'hfe;
      17'd46625: data = 8'hfe;
      17'd46626: data = 8'hfe;
      17'd46627: data = 8'hfd;
      17'd46628: data = 8'hfd;
      17'd46629: data = 8'hfd;
      17'd46630: data = 8'hfe;
      17'd46631: data = 8'h00;
      17'd46632: data = 8'hfe;
      17'd46633: data = 8'h00;
      17'd46634: data = 8'h00;
      17'd46635: data = 8'hfe;
      17'd46636: data = 8'hfe;
      17'd46637: data = 8'hfe;
      17'd46638: data = 8'hfd;
      17'd46639: data = 8'hfd;
      17'd46640: data = 8'hfe;
      17'd46641: data = 8'h00;
      17'd46642: data = 8'hfe;
      17'd46643: data = 8'hfe;
      17'd46644: data = 8'hfe;
      17'd46645: data = 8'h01;
      17'd46646: data = 8'h00;
      17'd46647: data = 8'hfe;
      17'd46648: data = 8'h00;
      17'd46649: data = 8'h00;
      17'd46650: data = 8'h00;
      17'd46651: data = 8'h00;
      17'd46652: data = 8'h00;
      17'd46653: data = 8'hfe;
      17'd46654: data = 8'hfe;
      17'd46655: data = 8'hfe;
      17'd46656: data = 8'hfd;
      17'd46657: data = 8'hfd;
      17'd46658: data = 8'hfe;
      17'd46659: data = 8'hfd;
      17'd46660: data = 8'h00;
      17'd46661: data = 8'h00;
      17'd46662: data = 8'h00;
      17'd46663: data = 8'h00;
      17'd46664: data = 8'hfe;
      17'd46665: data = 8'h00;
      17'd46666: data = 8'hfe;
      17'd46667: data = 8'hfe;
      17'd46668: data = 8'hfd;
      17'd46669: data = 8'hfd;
      17'd46670: data = 8'hfc;
      17'd46671: data = 8'hfd;
      17'd46672: data = 8'hfd;
      17'd46673: data = 8'hfd;
      17'd46674: data = 8'h00;
      17'd46675: data = 8'h00;
      17'd46676: data = 8'hfe;
      17'd46677: data = 8'h00;
      17'd46678: data = 8'h00;
      17'd46679: data = 8'h00;
      17'd46680: data = 8'h01;
      17'd46681: data = 8'h00;
      17'd46682: data = 8'h00;
      17'd46683: data = 8'h00;
      17'd46684: data = 8'hfd;
      17'd46685: data = 8'hfd;
      17'd46686: data = 8'hfe;
      17'd46687: data = 8'hfe;
      17'd46688: data = 8'hfe;
      17'd46689: data = 8'h00;
      17'd46690: data = 8'hfe;
      17'd46691: data = 8'h00;
      17'd46692: data = 8'h01;
      17'd46693: data = 8'h02;
      17'd46694: data = 8'h02;
      17'd46695: data = 8'h00;
      17'd46696: data = 8'hfe;
      17'd46697: data = 8'h00;
      17'd46698: data = 8'h01;
      17'd46699: data = 8'hfe;
      17'd46700: data = 8'hfe;
      17'd46701: data = 8'h00;
      17'd46702: data = 8'h00;
      17'd46703: data = 8'h01;
      17'd46704: data = 8'h00;
      17'd46705: data = 8'h00;
      17'd46706: data = 8'hfe;
      17'd46707: data = 8'h00;
      17'd46708: data = 8'h01;
      17'd46709: data = 8'h00;
      17'd46710: data = 8'h00;
      17'd46711: data = 8'hfe;
      17'd46712: data = 8'hfe;
      17'd46713: data = 8'h00;
      17'd46714: data = 8'h00;
      17'd46715: data = 8'h00;
      17'd46716: data = 8'hfd;
      17'd46717: data = 8'hfd;
      17'd46718: data = 8'hfe;
      17'd46719: data = 8'hfe;
      17'd46720: data = 8'hfe;
      17'd46721: data = 8'hfe;
      17'd46722: data = 8'h00;
      17'd46723: data = 8'h00;
      17'd46724: data = 8'h00;
      17'd46725: data = 8'h00;
      17'd46726: data = 8'h00;
      17'd46727: data = 8'h00;
      17'd46728: data = 8'hfe;
      17'd46729: data = 8'hfe;
      17'd46730: data = 8'h00;
      17'd46731: data = 8'h00;
      17'd46732: data = 8'hfe;
      17'd46733: data = 8'h00;
      17'd46734: data = 8'h00;
      17'd46735: data = 8'h01;
      17'd46736: data = 8'h00;
      17'd46737: data = 8'h00;
      17'd46738: data = 8'h01;
      17'd46739: data = 8'h00;
      17'd46740: data = 8'h00;
      17'd46741: data = 8'h00;
      17'd46742: data = 8'h00;
      17'd46743: data = 8'hfe;
      17'd46744: data = 8'hfe;
      17'd46745: data = 8'h00;
      17'd46746: data = 8'hfe;
      17'd46747: data = 8'hfe;
      17'd46748: data = 8'h00;
      17'd46749: data = 8'h00;
      17'd46750: data = 8'h00;
      17'd46751: data = 8'h01;
      17'd46752: data = 8'h00;
      17'd46753: data = 8'h00;
      17'd46754: data = 8'h01;
      17'd46755: data = 8'h01;
      17'd46756: data = 8'h00;
      17'd46757: data = 8'hfe;
      17'd46758: data = 8'hfe;
      17'd46759: data = 8'hfe;
      17'd46760: data = 8'hfe;
      17'd46761: data = 8'h00;
      17'd46762: data = 8'h00;
      17'd46763: data = 8'hfe;
      17'd46764: data = 8'hfe;
      17'd46765: data = 8'hfe;
      17'd46766: data = 8'hfd;
      17'd46767: data = 8'h00;
      17'd46768: data = 8'h01;
      17'd46769: data = 8'h00;
      17'd46770: data = 8'hfe;
      17'd46771: data = 8'h00;
      17'd46772: data = 8'h00;
      17'd46773: data = 8'hfe;
      17'd46774: data = 8'hfe;
      17'd46775: data = 8'hfe;
      17'd46776: data = 8'h00;
      17'd46777: data = 8'hfe;
      17'd46778: data = 8'h00;
      17'd46779: data = 8'h00;
      17'd46780: data = 8'hfe;
      17'd46781: data = 8'h00;
      17'd46782: data = 8'h01;
      17'd46783: data = 8'h00;
      17'd46784: data = 8'h00;
      17'd46785: data = 8'h00;
      17'd46786: data = 8'h00;
      17'd46787: data = 8'h00;
      17'd46788: data = 8'h00;
      17'd46789: data = 8'hfe;
      17'd46790: data = 8'hfd;
      17'd46791: data = 8'hfe;
      17'd46792: data = 8'hfe;
      17'd46793: data = 8'h00;
      17'd46794: data = 8'hfe;
      17'd46795: data = 8'hfe;
      17'd46796: data = 8'hfe;
      17'd46797: data = 8'h00;
      17'd46798: data = 8'h00;
      17'd46799: data = 8'h00;
      17'd46800: data = 8'hfe;
      17'd46801: data = 8'hfe;
      17'd46802: data = 8'h00;
      17'd46803: data = 8'hfe;
      17'd46804: data = 8'hfd;
      17'd46805: data = 8'hfe;
      17'd46806: data = 8'hfe;
      17'd46807: data = 8'hfe;
      17'd46808: data = 8'h00;
      17'd46809: data = 8'hfe;
      17'd46810: data = 8'hfd;
      17'd46811: data = 8'h00;
      17'd46812: data = 8'h00;
      17'd46813: data = 8'hfe;
      17'd46814: data = 8'hfe;
      17'd46815: data = 8'hfe;
      17'd46816: data = 8'hfe;
      17'd46817: data = 8'h00;
      17'd46818: data = 8'hfe;
      17'd46819: data = 8'hfe;
      17'd46820: data = 8'hfe;
      17'd46821: data = 8'hfe;
      17'd46822: data = 8'hfd;
      17'd46823: data = 8'hfe;
      17'd46824: data = 8'hfe;
      17'd46825: data = 8'hfe;
      17'd46826: data = 8'hfe;
      17'd46827: data = 8'hfe;
      17'd46828: data = 8'hfe;
      17'd46829: data = 8'hfe;
      17'd46830: data = 8'hfe;
      17'd46831: data = 8'h00;
      17'd46832: data = 8'hfe;
      17'd46833: data = 8'hfd;
      17'd46834: data = 8'hfe;
      17'd46835: data = 8'hfd;
      17'd46836: data = 8'hfe;
      17'd46837: data = 8'h00;
      17'd46838: data = 8'hfe;
      17'd46839: data = 8'hfe;
      17'd46840: data = 8'h00;
      17'd46841: data = 8'h00;
      17'd46842: data = 8'h00;
      17'd46843: data = 8'h00;
      17'd46844: data = 8'hfe;
      17'd46845: data = 8'h00;
      17'd46846: data = 8'h00;
      17'd46847: data = 8'h00;
      17'd46848: data = 8'h01;
      17'd46849: data = 8'h00;
      17'd46850: data = 8'hfe;
      17'd46851: data = 8'hfd;
      17'd46852: data = 8'hfe;
      17'd46853: data = 8'hfe;
      17'd46854: data = 8'h01;
      17'd46855: data = 8'h00;
      17'd46856: data = 8'hfe;
      17'd46857: data = 8'h00;
      17'd46858: data = 8'h00;
      17'd46859: data = 8'h01;
      17'd46860: data = 8'h02;
      17'd46861: data = 8'h01;
      17'd46862: data = 8'h00;
      17'd46863: data = 8'h00;
      17'd46864: data = 8'h01;
      17'd46865: data = 8'hfe;
      17'd46866: data = 8'hfe;
      17'd46867: data = 8'h00;
      17'd46868: data = 8'h00;
      17'd46869: data = 8'h00;
      17'd46870: data = 8'hfe;
      17'd46871: data = 8'h01;
      17'd46872: data = 8'h01;
      17'd46873: data = 8'h00;
      17'd46874: data = 8'h01;
      17'd46875: data = 8'h00;
      17'd46876: data = 8'h01;
      17'd46877: data = 8'h00;
      17'd46878: data = 8'h00;
      17'd46879: data = 8'hfd;
      17'd46880: data = 8'h00;
      17'd46881: data = 8'h00;
      17'd46882: data = 8'h00;
      17'd46883: data = 8'hfe;
      17'd46884: data = 8'hfd;
      17'd46885: data = 8'hfe;
      17'd46886: data = 8'h00;
      17'd46887: data = 8'h01;
      17'd46888: data = 8'h01;
      17'd46889: data = 8'h01;
      17'd46890: data = 8'h02;
      17'd46891: data = 8'h04;
      17'd46892: data = 8'h01;
      17'd46893: data = 8'h01;
      17'd46894: data = 8'h00;
      17'd46895: data = 8'h00;
      17'd46896: data = 8'hfe;
      17'd46897: data = 8'hfe;
      17'd46898: data = 8'hfe;
      17'd46899: data = 8'hfe;
      17'd46900: data = 8'hfe;
      17'd46901: data = 8'h00;
      17'd46902: data = 8'h01;
      17'd46903: data = 8'h00;
      17'd46904: data = 8'h01;
      17'd46905: data = 8'h02;
      17'd46906: data = 8'h01;
      17'd46907: data = 8'h01;
      17'd46908: data = 8'h01;
      17'd46909: data = 8'h01;
      17'd46910: data = 8'h00;
      17'd46911: data = 8'h00;
      17'd46912: data = 8'hfe;
      17'd46913: data = 8'hfe;
      17'd46914: data = 8'h00;
      17'd46915: data = 8'h00;
      17'd46916: data = 8'h00;
      17'd46917: data = 8'hfe;
      17'd46918: data = 8'hfe;
      17'd46919: data = 8'h00;
      17'd46920: data = 8'h01;
      17'd46921: data = 8'h01;
      17'd46922: data = 8'h00;
      17'd46923: data = 8'hfe;
      17'd46924: data = 8'hfe;
      17'd46925: data = 8'h00;
      17'd46926: data = 8'hfe;
      17'd46927: data = 8'hfe;
      17'd46928: data = 8'hfe;
      17'd46929: data = 8'hfd;
      17'd46930: data = 8'hfd;
      17'd46931: data = 8'hfd;
      17'd46932: data = 8'hfd;
      17'd46933: data = 8'hfd;
      17'd46934: data = 8'hfd;
      17'd46935: data = 8'hfd;
      17'd46936: data = 8'hfe;
      17'd46937: data = 8'h00;
      17'd46938: data = 8'h00;
      17'd46939: data = 8'h00;
      17'd46940: data = 8'h00;
      17'd46941: data = 8'h01;
      17'd46942: data = 8'h00;
      17'd46943: data = 8'h00;
      17'd46944: data = 8'h00;
      17'd46945: data = 8'hfe;
      17'd46946: data = 8'h00;
      17'd46947: data = 8'h00;
      17'd46948: data = 8'hfe;
      17'd46949: data = 8'h00;
      17'd46950: data = 8'h00;
      17'd46951: data = 8'h00;
      17'd46952: data = 8'h00;
      17'd46953: data = 8'h01;
      17'd46954: data = 8'h02;
      17'd46955: data = 8'h01;
      17'd46956: data = 8'h01;
      17'd46957: data = 8'hfe;
      17'd46958: data = 8'h00;
      17'd46959: data = 8'hfe;
      17'd46960: data = 8'hfe;
      17'd46961: data = 8'hfe;
      17'd46962: data = 8'hfe;
      17'd46963: data = 8'hfe;
      17'd46964: data = 8'hfe;
      17'd46965: data = 8'h00;
      17'd46966: data = 8'h01;
      17'd46967: data = 8'h01;
      17'd46968: data = 8'h01;
      17'd46969: data = 8'h01;
      17'd46970: data = 8'h01;
      17'd46971: data = 8'h01;
      17'd46972: data = 8'h01;
      17'd46973: data = 8'h00;
      17'd46974: data = 8'hfe;
      17'd46975: data = 8'hfe;
      17'd46976: data = 8'hfd;
      17'd46977: data = 8'hfe;
      17'd46978: data = 8'hfe;
      17'd46979: data = 8'h00;
      17'd46980: data = 8'h00;
      17'd46981: data = 8'h00;
      17'd46982: data = 8'h01;
      17'd46983: data = 8'h01;
      17'd46984: data = 8'h01;
      17'd46985: data = 8'h00;
      17'd46986: data = 8'h00;
      17'd46987: data = 8'h00;
      17'd46988: data = 8'h00;
      17'd46989: data = 8'h00;
      17'd46990: data = 8'hfe;
      17'd46991: data = 8'hfc;
      17'd46992: data = 8'hfe;
      17'd46993: data = 8'hfe;
      17'd46994: data = 8'hfe;
      17'd46995: data = 8'hfe;
      17'd46996: data = 8'hfe;
      17'd46997: data = 8'h00;
      17'd46998: data = 8'h00;
      17'd46999: data = 8'h02;
      17'd47000: data = 8'h01;
      17'd47001: data = 8'h01;
      17'd47002: data = 8'h01;
      17'd47003: data = 8'h00;
      17'd47004: data = 8'h00;
      17'd47005: data = 8'hfe;
      17'd47006: data = 8'hfe;
      17'd47007: data = 8'hfe;
      17'd47008: data = 8'h00;
      17'd47009: data = 8'h00;
      17'd47010: data = 8'h00;
      17'd47011: data = 8'h00;
      17'd47012: data = 8'h00;
      17'd47013: data = 8'h00;
      17'd47014: data = 8'h00;
      17'd47015: data = 8'h00;
      17'd47016: data = 8'h00;
      17'd47017: data = 8'h00;
      17'd47018: data = 8'h00;
      17'd47019: data = 8'hfe;
      17'd47020: data = 8'hfe;
      17'd47021: data = 8'hfe;
      17'd47022: data = 8'h00;
      17'd47023: data = 8'h00;
      17'd47024: data = 8'h00;
      17'd47025: data = 8'h01;
      17'd47026: data = 8'hfe;
      17'd47027: data = 8'hfe;
      17'd47028: data = 8'hfe;
      17'd47029: data = 8'hfe;
      17'd47030: data = 8'hfe;
      17'd47031: data = 8'hfe;
      17'd47032: data = 8'h00;
      17'd47033: data = 8'hfe;
      17'd47034: data = 8'h00;
      17'd47035: data = 8'hfe;
      17'd47036: data = 8'hfe;
      17'd47037: data = 8'h00;
      17'd47038: data = 8'h00;
      17'd47039: data = 8'h00;
      17'd47040: data = 8'h01;
      17'd47041: data = 8'h00;
      17'd47042: data = 8'hfe;
      17'd47043: data = 8'hfe;
      17'd47044: data = 8'hfe;
      17'd47045: data = 8'hfd;
      17'd47046: data = 8'hfd;
      17'd47047: data = 8'hfd;
      17'd47048: data = 8'h00;
      17'd47049: data = 8'h00;
      17'd47050: data = 8'h00;
      17'd47051: data = 8'h01;
      17'd47052: data = 8'h01;
      17'd47053: data = 8'h01;
      17'd47054: data = 8'h01;
      17'd47055: data = 8'h00;
      17'd47056: data = 8'hfe;
      17'd47057: data = 8'hfd;
      17'd47058: data = 8'hfd;
      17'd47059: data = 8'hfe;
      17'd47060: data = 8'hfd;
      17'd47061: data = 8'hfc;
      17'd47062: data = 8'hfc;
      17'd47063: data = 8'hfe;
      17'd47064: data = 8'h00;
      17'd47065: data = 8'hfe;
      17'd47066: data = 8'hfe;
      17'd47067: data = 8'hfe;
      17'd47068: data = 8'hfe;
      17'd47069: data = 8'hfe;
      17'd47070: data = 8'hfe;
      17'd47071: data = 8'hfd;
      17'd47072: data = 8'hfc;
      17'd47073: data = 8'hfc;
      17'd47074: data = 8'hfc;
      17'd47075: data = 8'hfc;
      17'd47076: data = 8'hfd;
      17'd47077: data = 8'hfe;
      17'd47078: data = 8'hfe;
      17'd47079: data = 8'h00;
      17'd47080: data = 8'hfe;
      17'd47081: data = 8'h00;
      17'd47082: data = 8'h01;
      17'd47083: data = 8'h01;
      17'd47084: data = 8'h00;
      17'd47085: data = 8'hfe;
      17'd47086: data = 8'hfe;
      17'd47087: data = 8'hfd;
      17'd47088: data = 8'hfd;
      17'd47089: data = 8'hfc;
      17'd47090: data = 8'hfd;
      17'd47091: data = 8'hfe;
      17'd47092: data = 8'hfd;
      17'd47093: data = 8'h00;
      17'd47094: data = 8'h01;
      17'd47095: data = 8'h02;
      17'd47096: data = 8'h02;
      17'd47097: data = 8'h01;
      17'd47098: data = 8'h02;
      17'd47099: data = 8'h01;
      17'd47100: data = 8'h00;
      17'd47101: data = 8'hfe;
      17'd47102: data = 8'hfc;
      17'd47103: data = 8'hfc;
      17'd47104: data = 8'hfd;
      17'd47105: data = 8'hfe;
      17'd47106: data = 8'hfd;
      17'd47107: data = 8'hfe;
      17'd47108: data = 8'h00;
      17'd47109: data = 8'h01;
      17'd47110: data = 8'h01;
      17'd47111: data = 8'h01;
      17'd47112: data = 8'h01;
      17'd47113: data = 8'h01;
      17'd47114: data = 8'h01;
      17'd47115: data = 8'h00;
      17'd47116: data = 8'h00;
      17'd47117: data = 8'hfd;
      17'd47118: data = 8'hfc;
      17'd47119: data = 8'hfd;
      17'd47120: data = 8'hfe;
      17'd47121: data = 8'h00;
      17'd47122: data = 8'h00;
      17'd47123: data = 8'h01;
      17'd47124: data = 8'h02;
      17'd47125: data = 8'h04;
      17'd47126: data = 8'h04;
      17'd47127: data = 8'h02;
      17'd47128: data = 8'h02;
      17'd47129: data = 8'h01;
      17'd47130: data = 8'h01;
      17'd47131: data = 8'h00;
      17'd47132: data = 8'hfe;
      17'd47133: data = 8'hfe;
      17'd47134: data = 8'h00;
      17'd47135: data = 8'hfe;
      17'd47136: data = 8'h00;
      17'd47137: data = 8'h01;
      17'd47138: data = 8'h01;
      17'd47139: data = 8'h02;
      17'd47140: data = 8'h02;
      17'd47141: data = 8'h02;
      17'd47142: data = 8'h04;
      17'd47143: data = 8'h02;
      17'd47144: data = 8'h00;
      17'd47145: data = 8'h01;
      17'd47146: data = 8'h01;
      17'd47147: data = 8'h00;
      17'd47148: data = 8'h00;
      17'd47149: data = 8'hfe;
      17'd47150: data = 8'h00;
      17'd47151: data = 8'h00;
      17'd47152: data = 8'h01;
      17'd47153: data = 8'h02;
      17'd47154: data = 8'h02;
      17'd47155: data = 8'h00;
      17'd47156: data = 8'h00;
      17'd47157: data = 8'h01;
      17'd47158: data = 8'h01;
      17'd47159: data = 8'h01;
      17'd47160: data = 8'h00;
      17'd47161: data = 8'h00;
      17'd47162: data = 8'hfd;
      17'd47163: data = 8'hfe;
      17'd47164: data = 8'hfe;
      17'd47165: data = 8'h00;
      17'd47166: data = 8'h00;
      17'd47167: data = 8'h01;
      17'd47168: data = 8'h01;
      17'd47169: data = 8'h01;
      17'd47170: data = 8'h02;
      17'd47171: data = 8'h01;
      17'd47172: data = 8'h00;
      17'd47173: data = 8'h00;
      17'd47174: data = 8'hfe;
      17'd47175: data = 8'h00;
      17'd47176: data = 8'hfe;
      17'd47177: data = 8'hfe;
      17'd47178: data = 8'hfe;
      17'd47179: data = 8'hfd;
      17'd47180: data = 8'h00;
      17'd47181: data = 8'h00;
      17'd47182: data = 8'h00;
      17'd47183: data = 8'h01;
      17'd47184: data = 8'h02;
      17'd47185: data = 8'h02;
      17'd47186: data = 8'h01;
      17'd47187: data = 8'hfe;
      17'd47188: data = 8'hfd;
      17'd47189: data = 8'hfd;
      17'd47190: data = 8'hfe;
      17'd47191: data = 8'hfd;
      17'd47192: data = 8'hfd;
      17'd47193: data = 8'hfe;
      17'd47194: data = 8'hfe;
      17'd47195: data = 8'h01;
      17'd47196: data = 8'h00;
      17'd47197: data = 8'h00;
      17'd47198: data = 8'h00;
      17'd47199: data = 8'h00;
      17'd47200: data = 8'h00;
      17'd47201: data = 8'hfd;
      17'd47202: data = 8'hfd;
      17'd47203: data = 8'hfd;
      17'd47204: data = 8'hfe;
      17'd47205: data = 8'hfe;
      17'd47206: data = 8'hfd;
      17'd47207: data = 8'hfe;
      17'd47208: data = 8'hfd;
      17'd47209: data = 8'hfe;
      17'd47210: data = 8'h00;
      17'd47211: data = 8'h00;
      17'd47212: data = 8'h00;
      17'd47213: data = 8'h00;
      17'd47214: data = 8'hfe;
      17'd47215: data = 8'h00;
      17'd47216: data = 8'h00;
      17'd47217: data = 8'hfe;
      17'd47218: data = 8'hfe;
      17'd47219: data = 8'hfd;
      17'd47220: data = 8'hfe;
      17'd47221: data = 8'hfe;
      17'd47222: data = 8'hfe;
      17'd47223: data = 8'hfe;
      17'd47224: data = 8'hfe;
      17'd47225: data = 8'h00;
      17'd47226: data = 8'h01;
      17'd47227: data = 8'h00;
      17'd47228: data = 8'h00;
      17'd47229: data = 8'h00;
      17'd47230: data = 8'hfd;
      17'd47231: data = 8'hfe;
      17'd47232: data = 8'h00;
      17'd47233: data = 8'hfe;
      17'd47234: data = 8'hfe;
      17'd47235: data = 8'hfd;
      17'd47236: data = 8'hfe;
      17'd47237: data = 8'h00;
      17'd47238: data = 8'h01;
      17'd47239: data = 8'h00;
      17'd47240: data = 8'h01;
      17'd47241: data = 8'h01;
      17'd47242: data = 8'h01;
      17'd47243: data = 8'h01;
      17'd47244: data = 8'hfe;
      17'd47245: data = 8'hfe;
      17'd47246: data = 8'hfe;
      17'd47247: data = 8'hfc;
      17'd47248: data = 8'hfa;
      17'd47249: data = 8'hfc;
      17'd47250: data = 8'hfd;
      17'd47251: data = 8'hfd;
      17'd47252: data = 8'hfe;
      17'd47253: data = 8'hfd;
      17'd47254: data = 8'hfe;
      17'd47255: data = 8'h01;
      17'd47256: data = 8'h00;
      17'd47257: data = 8'h00;
      17'd47258: data = 8'h01;
      17'd47259: data = 8'h00;
      17'd47260: data = 8'hfe;
      17'd47261: data = 8'hfd;
      17'd47262: data = 8'hfc;
      17'd47263: data = 8'hfd;
      17'd47264: data = 8'hfd;
      17'd47265: data = 8'hfd;
      17'd47266: data = 8'hfd;
      17'd47267: data = 8'hfd;
      17'd47268: data = 8'hfd;
      17'd47269: data = 8'h00;
      17'd47270: data = 8'h01;
      17'd47271: data = 8'h01;
      17'd47272: data = 8'h01;
      17'd47273: data = 8'h01;
      17'd47274: data = 8'h00;
      17'd47275: data = 8'hfe;
      17'd47276: data = 8'hfe;
      17'd47277: data = 8'hfd;
      17'd47278: data = 8'hfd;
      17'd47279: data = 8'hfe;
      17'd47280: data = 8'hfe;
      17'd47281: data = 8'hfd;
      17'd47282: data = 8'hfd;
      17'd47283: data = 8'hfd;
      17'd47284: data = 8'h00;
      17'd47285: data = 8'hfe;
      17'd47286: data = 8'h01;
      17'd47287: data = 8'h02;
      17'd47288: data = 8'h02;
      17'd47289: data = 8'h02;
      17'd47290: data = 8'h00;
      17'd47291: data = 8'h00;
      17'd47292: data = 8'hfe;
      17'd47293: data = 8'hfe;
      17'd47294: data = 8'hfd;
      17'd47295: data = 8'hfc;
      17'd47296: data = 8'hfd;
      17'd47297: data = 8'hfe;
      17'd47298: data = 8'hfe;
      17'd47299: data = 8'h00;
      17'd47300: data = 8'h00;
      17'd47301: data = 8'h01;
      17'd47302: data = 8'h02;
      17'd47303: data = 8'h01;
      17'd47304: data = 8'h00;
      17'd47305: data = 8'h00;
      17'd47306: data = 8'hfe;
      17'd47307: data = 8'hfe;
      17'd47308: data = 8'hfe;
      17'd47309: data = 8'hfd;
      17'd47310: data = 8'hfe;
      17'd47311: data = 8'hfd;
      17'd47312: data = 8'hfe;
      17'd47313: data = 8'hfe;
      17'd47314: data = 8'hfe;
      17'd47315: data = 8'h01;
      17'd47316: data = 8'h01;
      17'd47317: data = 8'h02;
      17'd47318: data = 8'h01;
      17'd47319: data = 8'h00;
      17'd47320: data = 8'hfe;
      17'd47321: data = 8'hfd;
      17'd47322: data = 8'hfd;
      17'd47323: data = 8'hfd;
      17'd47324: data = 8'hfc;
      17'd47325: data = 8'hfc;
      17'd47326: data = 8'hfd;
      17'd47327: data = 8'hfd;
      17'd47328: data = 8'hfe;
      17'd47329: data = 8'hfe;
      17'd47330: data = 8'h00;
      17'd47331: data = 8'h01;
      17'd47332: data = 8'h01;
      17'd47333: data = 8'h00;
      17'd47334: data = 8'hfe;
      17'd47335: data = 8'h00;
      17'd47336: data = 8'h00;
      17'd47337: data = 8'hfe;
      17'd47338: data = 8'hfe;
      17'd47339: data = 8'hfd;
      17'd47340: data = 8'hfd;
      17'd47341: data = 8'hfe;
      17'd47342: data = 8'hfe;
      17'd47343: data = 8'hfe;
      17'd47344: data = 8'h00;
      17'd47345: data = 8'h01;
      17'd47346: data = 8'h02;
      17'd47347: data = 8'h02;
      17'd47348: data = 8'h02;
      17'd47349: data = 8'h01;
      17'd47350: data = 8'h01;
      17'd47351: data = 8'h00;
      17'd47352: data = 8'h00;
      17'd47353: data = 8'h00;
      17'd47354: data = 8'hfe;
      17'd47355: data = 8'h00;
      17'd47356: data = 8'h00;
      17'd47357: data = 8'h00;
      17'd47358: data = 8'h00;
      17'd47359: data = 8'h01;
      17'd47360: data = 8'h01;
      17'd47361: data = 8'h02;
      17'd47362: data = 8'h01;
      17'd47363: data = 8'h01;
      17'd47364: data = 8'h01;
      17'd47365: data = 8'h01;
      17'd47366: data = 8'h01;
      17'd47367: data = 8'h01;
      17'd47368: data = 8'h00;
      17'd47369: data = 8'h00;
      17'd47370: data = 8'h01;
      17'd47371: data = 8'h01;
      17'd47372: data = 8'h00;
      17'd47373: data = 8'h01;
      17'd47374: data = 8'h01;
      17'd47375: data = 8'h02;
      17'd47376: data = 8'h01;
      17'd47377: data = 8'h02;
      17'd47378: data = 8'h01;
      17'd47379: data = 8'h00;
      17'd47380: data = 8'h00;
      17'd47381: data = 8'h00;
      17'd47382: data = 8'h00;
      17'd47383: data = 8'h01;
      17'd47384: data = 8'h01;
      17'd47385: data = 8'h00;
      17'd47386: data = 8'h02;
      17'd47387: data = 8'h02;
      17'd47388: data = 8'h02;
      17'd47389: data = 8'h04;
      17'd47390: data = 8'h04;
      17'd47391: data = 8'h04;
      17'd47392: data = 8'h02;
      17'd47393: data = 8'h02;
      17'd47394: data = 8'h01;
      17'd47395: data = 8'h00;
      17'd47396: data = 8'hfe;
      17'd47397: data = 8'h00;
      17'd47398: data = 8'h01;
      17'd47399: data = 8'h00;
      17'd47400: data = 8'h01;
      17'd47401: data = 8'h02;
      17'd47402: data = 8'h01;
      17'd47403: data = 8'h02;
      17'd47404: data = 8'h04;
      17'd47405: data = 8'h02;
      17'd47406: data = 8'h01;
      17'd47407: data = 8'h00;
      17'd47408: data = 8'h00;
      17'd47409: data = 8'h01;
      17'd47410: data = 8'hfe;
      17'd47411: data = 8'hfe;
      17'd47412: data = 8'hfe;
      17'd47413: data = 8'h00;
      17'd47414: data = 8'h00;
      17'd47415: data = 8'hfe;
      17'd47416: data = 8'hfe;
      17'd47417: data = 8'h00;
      17'd47418: data = 8'h02;
      17'd47419: data = 8'h01;
      17'd47420: data = 8'h01;
      17'd47421: data = 8'h01;
      17'd47422: data = 8'h01;
      17'd47423: data = 8'h01;
      17'd47424: data = 8'hfd;
      17'd47425: data = 8'hfc;
      17'd47426: data = 8'hfe;
      17'd47427: data = 8'hfd;
      17'd47428: data = 8'hfd;
      17'd47429: data = 8'hfe;
      17'd47430: data = 8'hfe;
      17'd47431: data = 8'hfe;
      17'd47432: data = 8'h00;
      17'd47433: data = 8'h00;
      17'd47434: data = 8'h01;
      17'd47435: data = 8'h01;
      17'd47436: data = 8'h00;
      17'd47437: data = 8'h01;
      17'd47438: data = 8'h00;
      17'd47439: data = 8'hfe;
      17'd47440: data = 8'hfe;
      17'd47441: data = 8'hfe;
      17'd47442: data = 8'h00;
      17'd47443: data = 8'hfe;
      17'd47444: data = 8'hfe;
      17'd47445: data = 8'hfe;
      17'd47446: data = 8'hfe;
      17'd47447: data = 8'hfe;
      17'd47448: data = 8'hfe;
      17'd47449: data = 8'hfe;
      17'd47450: data = 8'h00;
      17'd47451: data = 8'h00;
      17'd47452: data = 8'h00;
      17'd47453: data = 8'h00;
      17'd47454: data = 8'h00;
      17'd47455: data = 8'h00;
      17'd47456: data = 8'hfe;
      17'd47457: data = 8'hfe;
      17'd47458: data = 8'hfd;
      17'd47459: data = 8'hfc;
      17'd47460: data = 8'hfd;
      17'd47461: data = 8'hfd;
      17'd47462: data = 8'hfd;
      17'd47463: data = 8'hfe;
      17'd47464: data = 8'hfd;
      17'd47465: data = 8'h00;
      17'd47466: data = 8'h00;
      17'd47467: data = 8'h00;
      17'd47468: data = 8'h00;
      17'd47469: data = 8'hfe;
      17'd47470: data = 8'h00;
      17'd47471: data = 8'hfe;
      17'd47472: data = 8'hfd;
      17'd47473: data = 8'hfe;
      17'd47474: data = 8'hfe;
      17'd47475: data = 8'h00;
      17'd47476: data = 8'hfd;
      17'd47477: data = 8'hfd;
      17'd47478: data = 8'hfe;
      17'd47479: data = 8'h00;
      17'd47480: data = 8'h01;
      17'd47481: data = 8'h01;
      17'd47482: data = 8'h01;
      17'd47483: data = 8'h01;
      17'd47484: data = 8'h00;
      17'd47485: data = 8'h00;
      17'd47486: data = 8'h00;
      17'd47487: data = 8'hfe;
      17'd47488: data = 8'hfe;
      17'd47489: data = 8'hfe;
      17'd47490: data = 8'hfd;
      17'd47491: data = 8'hfe;
      17'd47492: data = 8'hfe;
      17'd47493: data = 8'h00;
      17'd47494: data = 8'hfe;
      17'd47495: data = 8'hfe;
      17'd47496: data = 8'h00;
      17'd47497: data = 8'hfe;
      17'd47498: data = 8'hfe;
      17'd47499: data = 8'h01;
      17'd47500: data = 8'h00;
      17'd47501: data = 8'hfd;
      17'd47502: data = 8'hfe;
      17'd47503: data = 8'hfd;
      17'd47504: data = 8'hfc;
      17'd47505: data = 8'hfc;
      17'd47506: data = 8'hfc;
      17'd47507: data = 8'hfd;
      17'd47508: data = 8'hfe;
      17'd47509: data = 8'h00;
      17'd47510: data = 8'hfd;
      17'd47511: data = 8'hfe;
      17'd47512: data = 8'h01;
      17'd47513: data = 8'hfe;
      17'd47514: data = 8'hfe;
      17'd47515: data = 8'hfe;
      17'd47516: data = 8'hfe;
      17'd47517: data = 8'h00;
      17'd47518: data = 8'hfe;
      17'd47519: data = 8'hfe;
      17'd47520: data = 8'hfd;
      17'd47521: data = 8'hfd;
      17'd47522: data = 8'hfe;
      17'd47523: data = 8'hfe;
      17'd47524: data = 8'h00;
      17'd47525: data = 8'h00;
      17'd47526: data = 8'h00;
      17'd47527: data = 8'h00;
      17'd47528: data = 8'h01;
      17'd47529: data = 8'h00;
      17'd47530: data = 8'h00;
      17'd47531: data = 8'hfe;
      17'd47532: data = 8'hfe;
      17'd47533: data = 8'h00;
      17'd47534: data = 8'hfe;
      17'd47535: data = 8'hfc;
      17'd47536: data = 8'hfe;
      17'd47537: data = 8'h00;
      17'd47538: data = 8'hfe;
      17'd47539: data = 8'h01;
      17'd47540: data = 8'h01;
      17'd47541: data = 8'h00;
      17'd47542: data = 8'h00;
      17'd47543: data = 8'h01;
      17'd47544: data = 8'hfe;
      17'd47545: data = 8'h00;
      17'd47546: data = 8'h00;
      17'd47547: data = 8'hfe;
      17'd47548: data = 8'hfe;
      17'd47549: data = 8'h00;
      17'd47550: data = 8'hfe;
      17'd47551: data = 8'hfe;
      17'd47552: data = 8'hfe;
      17'd47553: data = 8'hfe;
      17'd47554: data = 8'hfd;
      17'd47555: data = 8'hfe;
      17'd47556: data = 8'h00;
      17'd47557: data = 8'hfe;
      17'd47558: data = 8'hfe;
      17'd47559: data = 8'h00;
      17'd47560: data = 8'hfe;
      17'd47561: data = 8'hfe;
      17'd47562: data = 8'hfd;
      17'd47563: data = 8'hfe;
      17'd47564: data = 8'hfe;
      17'd47565: data = 8'hfd;
      17'd47566: data = 8'hfe;
      17'd47567: data = 8'hfe;
      17'd47568: data = 8'hfe;
      17'd47569: data = 8'h00;
      17'd47570: data = 8'h00;
      17'd47571: data = 8'hfe;
      17'd47572: data = 8'hfe;
      17'd47573: data = 8'h01;
      17'd47574: data = 8'h00;
      17'd47575: data = 8'hfd;
      17'd47576: data = 8'hfe;
      17'd47577: data = 8'hfe;
      17'd47578: data = 8'hfe;
      17'd47579: data = 8'hfe;
      17'd47580: data = 8'h00;
      17'd47581: data = 8'hfe;
      17'd47582: data = 8'h00;
      17'd47583: data = 8'hfe;
      17'd47584: data = 8'hfe;
      17'd47585: data = 8'hfe;
      17'd47586: data = 8'hfe;
      17'd47587: data = 8'h00;
      17'd47588: data = 8'hfe;
      17'd47589: data = 8'hfe;
      17'd47590: data = 8'h00;
      17'd47591: data = 8'hfe;
      17'd47592: data = 8'hfd;
      17'd47593: data = 8'hfd;
      17'd47594: data = 8'hfe;
      17'd47595: data = 8'hfe;
      17'd47596: data = 8'hfd;
      17'd47597: data = 8'hfd;
      17'd47598: data = 8'hfd;
      17'd47599: data = 8'hfd;
      17'd47600: data = 8'hfe;
      17'd47601: data = 8'h00;
      17'd47602: data = 8'hfe;
      17'd47603: data = 8'h00;
      17'd47604: data = 8'hfe;
      17'd47605: data = 8'hfd;
      17'd47606: data = 8'hfe;
      17'd47607: data = 8'hfe;
      17'd47608: data = 8'hfe;
      17'd47609: data = 8'hfd;
      17'd47610: data = 8'h00;
      17'd47611: data = 8'h00;
      17'd47612: data = 8'hfe;
      17'd47613: data = 8'hfe;
      17'd47614: data = 8'hfe;
      17'd47615: data = 8'hfe;
      17'd47616: data = 8'hfe;
      17'd47617: data = 8'h01;
      17'd47618: data = 8'h00;
      17'd47619: data = 8'hfe;
      17'd47620: data = 8'hfe;
      17'd47621: data = 8'h00;
      17'd47622: data = 8'h00;
      17'd47623: data = 8'hfe;
      17'd47624: data = 8'hfe;
      17'd47625: data = 8'hfe;
      17'd47626: data = 8'h00;
      17'd47627: data = 8'hfe;
      17'd47628: data = 8'hfe;
      17'd47629: data = 8'hfe;
      17'd47630: data = 8'hfd;
      17'd47631: data = 8'h00;
      17'd47632: data = 8'h01;
      17'd47633: data = 8'h00;
      17'd47634: data = 8'h00;
      17'd47635: data = 8'h00;
      17'd47636: data = 8'h00;
      17'd47637: data = 8'h00;
      17'd47638: data = 8'hfe;
      17'd47639: data = 8'h00;
      17'd47640: data = 8'h00;
      17'd47641: data = 8'hfe;
      17'd47642: data = 8'hfe;
      17'd47643: data = 8'hfd;
      17'd47644: data = 8'hfe;
      17'd47645: data = 8'hfe;
      17'd47646: data = 8'h00;
      17'd47647: data = 8'hfe;
      17'd47648: data = 8'hfe;
      17'd47649: data = 8'hfe;
      17'd47650: data = 8'h00;
      17'd47651: data = 8'h01;
      17'd47652: data = 8'h00;
      17'd47653: data = 8'h01;
      17'd47654: data = 8'h00;
      17'd47655: data = 8'h00;
      17'd47656: data = 8'h00;
      17'd47657: data = 8'hfe;
      17'd47658: data = 8'h01;
      17'd47659: data = 8'h01;
      17'd47660: data = 8'h00;
      17'd47661: data = 8'h00;
      17'd47662: data = 8'h00;
      17'd47663: data = 8'h00;
      17'd47664: data = 8'hfe;
      17'd47665: data = 8'h01;
      17'd47666: data = 8'h00;
      17'd47667: data = 8'hfe;
      17'd47668: data = 8'hfe;
      17'd47669: data = 8'h00;
      17'd47670: data = 8'h00;
      17'd47671: data = 8'h00;
      17'd47672: data = 8'h00;
      17'd47673: data = 8'h00;
      17'd47674: data = 8'h00;
      17'd47675: data = 8'h00;
      17'd47676: data = 8'h00;
      17'd47677: data = 8'hfe;
      17'd47678: data = 8'hfe;
      17'd47679: data = 8'h00;
      17'd47680: data = 8'h01;
      17'd47681: data = 8'h00;
      17'd47682: data = 8'hfe;
      17'd47683: data = 8'hfe;
      17'd47684: data = 8'h00;
      17'd47685: data = 8'h00;
      17'd47686: data = 8'h00;
      17'd47687: data = 8'hfe;
      17'd47688: data = 8'hfe;
      17'd47689: data = 8'hfe;
      17'd47690: data = 8'h00;
      17'd47691: data = 8'h00;
      17'd47692: data = 8'hfe;
      17'd47693: data = 8'hfe;
      17'd47694: data = 8'h01;
      17'd47695: data = 8'h01;
      17'd47696: data = 8'h01;
      17'd47697: data = 8'h00;
      17'd47698: data = 8'h00;
      17'd47699: data = 8'hfe;
      17'd47700: data = 8'h00;
      17'd47701: data = 8'h00;
      17'd47702: data = 8'hfe;
      17'd47703: data = 8'h00;
      17'd47704: data = 8'hfe;
      17'd47705: data = 8'hfd;
      17'd47706: data = 8'hfe;
      17'd47707: data = 8'h00;
      17'd47708: data = 8'hfe;
      17'd47709: data = 8'hfe;
      17'd47710: data = 8'h00;
      17'd47711: data = 8'hfe;
      17'd47712: data = 8'hfe;
      17'd47713: data = 8'hfe;
      17'd47714: data = 8'h00;
      17'd47715: data = 8'h00;
      17'd47716: data = 8'h01;
      17'd47717: data = 8'h00;
      17'd47718: data = 8'h00;
      17'd47719: data = 8'h00;
      17'd47720: data = 8'h00;
      17'd47721: data = 8'h00;
      17'd47722: data = 8'h00;
      17'd47723: data = 8'hfe;
      17'd47724: data = 8'h00;
      17'd47725: data = 8'hfe;
      17'd47726: data = 8'h00;
      17'd47727: data = 8'h00;
      17'd47728: data = 8'h00;
      17'd47729: data = 8'h00;
      17'd47730: data = 8'h00;
      17'd47731: data = 8'hfe;
      17'd47732: data = 8'h00;
      17'd47733: data = 8'h00;
      17'd47734: data = 8'hfe;
      17'd47735: data = 8'hfe;
      17'd47736: data = 8'h00;
      17'd47737: data = 8'hfe;
      17'd47738: data = 8'hfe;
      17'd47739: data = 8'hfe;
      17'd47740: data = 8'hfd;
      17'd47741: data = 8'hfd;
      17'd47742: data = 8'hfe;
      17'd47743: data = 8'hfe;
      17'd47744: data = 8'h00;
      17'd47745: data = 8'h00;
      17'd47746: data = 8'hfe;
      17'd47747: data = 8'h00;
      17'd47748: data = 8'h00;
      17'd47749: data = 8'h00;
      17'd47750: data = 8'hfe;
      17'd47751: data = 8'h01;
      17'd47752: data = 8'h00;
      17'd47753: data = 8'hfe;
      17'd47754: data = 8'h00;
      17'd47755: data = 8'h00;
      17'd47756: data = 8'h00;
      17'd47757: data = 8'hfe;
      17'd47758: data = 8'hfe;
      17'd47759: data = 8'h00;
      17'd47760: data = 8'h00;
      17'd47761: data = 8'h00;
      17'd47762: data = 8'hfe;
      17'd47763: data = 8'hfe;
      17'd47764: data = 8'hfe;
      17'd47765: data = 8'hfe;
      17'd47766: data = 8'h00;
      17'd47767: data = 8'hfe;
      17'd47768: data = 8'hfe;
      17'd47769: data = 8'hfe;
      17'd47770: data = 8'hfe;
      17'd47771: data = 8'hfe;
      17'd47772: data = 8'hfe;
      17'd47773: data = 8'h00;
      17'd47774: data = 8'h00;
      17'd47775: data = 8'hfe;
      17'd47776: data = 8'hfd;
      17'd47777: data = 8'hfe;
      17'd47778: data = 8'hfe;
      17'd47779: data = 8'hfe;
      17'd47780: data = 8'hfe;
      17'd47781: data = 8'hfe;
      17'd47782: data = 8'hfe;
      17'd47783: data = 8'h00;
      17'd47784: data = 8'h00;
      17'd47785: data = 8'hfe;
      17'd47786: data = 8'h00;
      17'd47787: data = 8'hfe;
      17'd47788: data = 8'h00;
      17'd47789: data = 8'h01;
      17'd47790: data = 8'h00;
      17'd47791: data = 8'h00;
      17'd47792: data = 8'h01;
      17'd47793: data = 8'h00;
      17'd47794: data = 8'hfe;
      17'd47795: data = 8'h01;
      17'd47796: data = 8'h00;
      17'd47797: data = 8'h00;
      17'd47798: data = 8'h00;
      17'd47799: data = 8'h00;
      17'd47800: data = 8'h00;
      17'd47801: data = 8'h00;
      17'd47802: data = 8'hfe;
      17'd47803: data = 8'hfe;
      17'd47804: data = 8'hfe;
      17'd47805: data = 8'h00;
      17'd47806: data = 8'h00;
      17'd47807: data = 8'h00;
      17'd47808: data = 8'h00;
      17'd47809: data = 8'hfe;
      17'd47810: data = 8'h00;
      17'd47811: data = 8'hfe;
      17'd47812: data = 8'hfe;
      17'd47813: data = 8'hfe;
      17'd47814: data = 8'hfe;
      17'd47815: data = 8'h00;
      17'd47816: data = 8'h00;
      17'd47817: data = 8'hfe;
      17'd47818: data = 8'hfe;
      17'd47819: data = 8'h00;
      17'd47820: data = 8'h00;
      17'd47821: data = 8'h00;
      17'd47822: data = 8'h00;
      17'd47823: data = 8'h00;
      17'd47824: data = 8'h00;
      17'd47825: data = 8'h00;
      17'd47826: data = 8'h00;
      17'd47827: data = 8'h00;
      17'd47828: data = 8'hfe;
      17'd47829: data = 8'hfe;
      17'd47830: data = 8'h00;
      17'd47831: data = 8'hfe;
      17'd47832: data = 8'hfe;
      17'd47833: data = 8'h00;
      17'd47834: data = 8'h00;
      17'd47835: data = 8'h00;
      17'd47836: data = 8'h01;
      17'd47837: data = 8'h00;
      17'd47838: data = 8'h00;
      17'd47839: data = 8'h00;
      17'd47840: data = 8'hfe;
      17'd47841: data = 8'h00;
      17'd47842: data = 8'hfe;
      17'd47843: data = 8'hfe;
      17'd47844: data = 8'h00;
      17'd47845: data = 8'h01;
      17'd47846: data = 8'hfe;
      17'd47847: data = 8'h00;
      17'd47848: data = 8'h00;
      17'd47849: data = 8'hfe;
      17'd47850: data = 8'hfe;
      17'd47851: data = 8'hfe;
      17'd47852: data = 8'hfd;
      17'd47853: data = 8'hfe;
      17'd47854: data = 8'hfe;
      17'd47855: data = 8'hfd;
      17'd47856: data = 8'hfe;
      17'd47857: data = 8'hfe;
      17'd47858: data = 8'h01;
      17'd47859: data = 8'h00;
      17'd47860: data = 8'hfe;
      17'd47861: data = 8'h00;
      17'd47862: data = 8'h00;
      17'd47863: data = 8'h00;
      17'd47864: data = 8'h00;
      17'd47865: data = 8'h00;
      17'd47866: data = 8'h00;
      17'd47867: data = 8'hfe;
      17'd47868: data = 8'hfe;
      17'd47869: data = 8'hfe;
      17'd47870: data = 8'hfe;
      17'd47871: data = 8'hfe;
      17'd47872: data = 8'hfe;
      17'd47873: data = 8'h00;
      17'd47874: data = 8'h00;
      17'd47875: data = 8'h00;
      17'd47876: data = 8'h01;
      17'd47877: data = 8'h00;
      17'd47878: data = 8'h00;
      17'd47879: data = 8'h00;
      17'd47880: data = 8'h00;
      17'd47881: data = 8'h00;
      17'd47882: data = 8'h00;
      17'd47883: data = 8'h00;
      17'd47884: data = 8'hfe;
      17'd47885: data = 8'hfd;
      17'd47886: data = 8'hfd;
      17'd47887: data = 8'hfe;
      17'd47888: data = 8'hfe;
      17'd47889: data = 8'hfe;
      17'd47890: data = 8'hfe;
      17'd47891: data = 8'hfe;
      17'd47892: data = 8'h00;
      17'd47893: data = 8'hfe;
      17'd47894: data = 8'h00;
      17'd47895: data = 8'hfe;
      17'd47896: data = 8'hfe;
      17'd47897: data = 8'h00;
      17'd47898: data = 8'hfe;
      17'd47899: data = 8'hfe;
      17'd47900: data = 8'hfe;
      17'd47901: data = 8'hfe;
      17'd47902: data = 8'hfd;
      17'd47903: data = 8'hfd;
      17'd47904: data = 8'hfe;
      17'd47905: data = 8'hfe;
      17'd47906: data = 8'h00;
      17'd47907: data = 8'h00;
      17'd47908: data = 8'hfe;
      17'd47909: data = 8'h00;
      17'd47910: data = 8'h01;
      17'd47911: data = 8'h00;
      17'd47912: data = 8'hfe;
      17'd47913: data = 8'hfe;
      17'd47914: data = 8'h00;
      17'd47915: data = 8'hfe;
      17'd47916: data = 8'hfe;
      17'd47917: data = 8'hfe;
      17'd47918: data = 8'hfe;
      17'd47919: data = 8'h00;
      17'd47920: data = 8'h00;
      17'd47921: data = 8'h00;
      17'd47922: data = 8'hfe;
      17'd47923: data = 8'hfe;
      17'd47924: data = 8'h00;
      17'd47925: data = 8'hfe;
      17'd47926: data = 8'h00;
      17'd47927: data = 8'hfe;
      17'd47928: data = 8'hfe;
      17'd47929: data = 8'h00;
      17'd47930: data = 8'h00;
      17'd47931: data = 8'h00;
      17'd47932: data = 8'hfe;
      17'd47933: data = 8'hfe;
      17'd47934: data = 8'h00;
      17'd47935: data = 8'h00;
      17'd47936: data = 8'hfe;
      17'd47937: data = 8'h01;
      17'd47938: data = 8'h00;
      17'd47939: data = 8'h00;
      17'd47940: data = 8'h00;
      17'd47941: data = 8'h00;
      17'd47942: data = 8'hfe;
      17'd47943: data = 8'h00;
      17'd47944: data = 8'h01;
      17'd47945: data = 8'hfe;
      17'd47946: data = 8'h00;
      17'd47947: data = 8'h00;
      17'd47948: data = 8'h00;
      17'd47949: data = 8'hfd;
      17'd47950: data = 8'h00;
      17'd47951: data = 8'h00;
      17'd47952: data = 8'h00;
      17'd47953: data = 8'h01;
      17'd47954: data = 8'h00;
      17'd47955: data = 8'h00;
      17'd47956: data = 8'h00;
      17'd47957: data = 8'h00;
      17'd47958: data = 8'h00;
      17'd47959: data = 8'h00;
      17'd47960: data = 8'h00;
      17'd47961: data = 8'h00;
      17'd47962: data = 8'h00;
      17'd47963: data = 8'h00;
      17'd47964: data = 8'h00;
      17'd47965: data = 8'hfe;
      17'd47966: data = 8'h00;
      17'd47967: data = 8'h00;
      17'd47968: data = 8'h00;
      17'd47969: data = 8'h01;
      17'd47970: data = 8'h01;
      17'd47971: data = 8'h01;
      17'd47972: data = 8'h01;
      17'd47973: data = 8'h00;
      17'd47974: data = 8'h00;
      17'd47975: data = 8'h00;
      17'd47976: data = 8'h00;
      17'd47977: data = 8'h01;
      17'd47978: data = 8'h00;
      17'd47979: data = 8'h00;
      17'd47980: data = 8'h00;
      17'd47981: data = 8'h00;
      17'd47982: data = 8'hfe;
      17'd47983: data = 8'h01;
      17'd47984: data = 8'h00;
      17'd47985: data = 8'hfe;
      17'd47986: data = 8'h00;
      17'd47987: data = 8'h00;
      17'd47988: data = 8'h00;
      17'd47989: data = 8'hfe;
      17'd47990: data = 8'hfc;
      17'd47991: data = 8'h00;
      17'd47992: data = 8'h00;
      17'd47993: data = 8'hfe;
      17'd47994: data = 8'hfe;
      17'd47995: data = 8'hfe;
      17'd47996: data = 8'h00;
      17'd47997: data = 8'hfe;
      17'd47998: data = 8'hfd;
      17'd47999: data = 8'hfd;
      17'd48000: data = 8'hfd;
      17'd48001: data = 8'hfe;
      17'd48002: data = 8'hfe;
      17'd48003: data = 8'hfe;
      17'd48004: data = 8'hfd;
      17'd48005: data = 8'hfe;
      17'd48006: data = 8'h00;
      17'd48007: data = 8'hfe;
      17'd48008: data = 8'hfe;
      17'd48009: data = 8'hfe;
      17'd48010: data = 8'hfd;
      17'd48011: data = 8'hfe;
      17'd48012: data = 8'h00;
      17'd48013: data = 8'hfe;
      17'd48014: data = 8'hfe;
      17'd48015: data = 8'hfe;
      17'd48016: data = 8'hfe;
      17'd48017: data = 8'hfe;
      17'd48018: data = 8'hfe;
      17'd48019: data = 8'hfe;
      17'd48020: data = 8'hfe;
      17'd48021: data = 8'h00;
      17'd48022: data = 8'h00;
      17'd48023: data = 8'hfe;
      17'd48024: data = 8'hfd;
      17'd48025: data = 8'hfe;
      17'd48026: data = 8'h00;
      17'd48027: data = 8'hfd;
      17'd48028: data = 8'h00;
      17'd48029: data = 8'hfe;
      17'd48030: data = 8'hfe;
      17'd48031: data = 8'hfe;
      17'd48032: data = 8'hfe;
      17'd48033: data = 8'hfe;
      17'd48034: data = 8'hfe;
      17'd48035: data = 8'h00;
      17'd48036: data = 8'hfe;
      17'd48037: data = 8'h00;
      17'd48038: data = 8'hfe;
      17'd48039: data = 8'h00;
      17'd48040: data = 8'hfe;
      17'd48041: data = 8'hfd;
      17'd48042: data = 8'hfe;
      17'd48043: data = 8'hfe;
      17'd48044: data = 8'h00;
      17'd48045: data = 8'hfe;
      17'd48046: data = 8'h00;
      17'd48047: data = 8'hfe;
      17'd48048: data = 8'hfe;
      17'd48049: data = 8'h00;
      17'd48050: data = 8'h01;
      17'd48051: data = 8'h01;
      17'd48052: data = 8'h01;
      17'd48053: data = 8'h01;
      17'd48054: data = 8'h00;
      17'd48055: data = 8'h00;
      17'd48056: data = 8'h00;
      17'd48057: data = 8'h00;
      17'd48058: data = 8'h00;
      17'd48059: data = 8'h00;
      17'd48060: data = 8'h00;
      17'd48061: data = 8'h00;
      17'd48062: data = 8'h02;
      17'd48063: data = 8'h01;
      17'd48064: data = 8'h01;
      17'd48065: data = 8'h01;
      17'd48066: data = 8'h00;
      17'd48067: data = 8'h00;
      17'd48068: data = 8'h00;
      17'd48069: data = 8'h01;
      17'd48070: data = 8'h00;
      17'd48071: data = 8'h00;
      17'd48072: data = 8'h00;
      17'd48073: data = 8'h01;
      17'd48074: data = 8'h00;
      17'd48075: data = 8'h00;
      17'd48076: data = 8'h00;
      17'd48077: data = 8'hfe;
      17'd48078: data = 8'hfe;
      17'd48079: data = 8'hfe;
      17'd48080: data = 8'h00;
      17'd48081: data = 8'h01;
      17'd48082: data = 8'h00;
      17'd48083: data = 8'hfe;
      17'd48084: data = 8'h01;
      17'd48085: data = 8'h01;
      17'd48086: data = 8'hfe;
      17'd48087: data = 8'h00;
      17'd48088: data = 8'h01;
      17'd48089: data = 8'h01;
      17'd48090: data = 8'h00;
      17'd48091: data = 8'h01;
      17'd48092: data = 8'h00;
      17'd48093: data = 8'h01;
      17'd48094: data = 8'h00;
      17'd48095: data = 8'hfe;
      17'd48096: data = 8'h00;
      17'd48097: data = 8'h00;
      17'd48098: data = 8'hfe;
      17'd48099: data = 8'hfd;
      17'd48100: data = 8'hfe;
      17'd48101: data = 8'hfe;
      17'd48102: data = 8'hfe;
      17'd48103: data = 8'h00;
      17'd48104: data = 8'h00;
      17'd48105: data = 8'h00;
      17'd48106: data = 8'h01;
      17'd48107: data = 8'h00;
      17'd48108: data = 8'h00;
      17'd48109: data = 8'h00;
      17'd48110: data = 8'hfe;
      17'd48111: data = 8'hfd;
      17'd48112: data = 8'hfd;
      17'd48113: data = 8'hfd;
      17'd48114: data = 8'hfd;
      17'd48115: data = 8'hfe;
      17'd48116: data = 8'hfd;
      17'd48117: data = 8'hfe;
      17'd48118: data = 8'hfe;
      17'd48119: data = 8'h00;
      17'd48120: data = 8'h00;
      17'd48121: data = 8'h00;
      17'd48122: data = 8'h00;
      17'd48123: data = 8'h00;
      17'd48124: data = 8'h00;
      17'd48125: data = 8'hfd;
      17'd48126: data = 8'hfd;
      17'd48127: data = 8'hfd;
      17'd48128: data = 8'hfd;
      17'd48129: data = 8'hfc;
      17'd48130: data = 8'hfd;
      17'd48131: data = 8'hfe;
      17'd48132: data = 8'hfe;
      17'd48133: data = 8'h00;
      17'd48134: data = 8'h00;
      17'd48135: data = 8'h00;
      17'd48136: data = 8'h00;
      17'd48137: data = 8'h01;
      17'd48138: data = 8'h00;
      17'd48139: data = 8'h00;
      17'd48140: data = 8'hfd;
      17'd48141: data = 8'hfd;
      17'd48142: data = 8'hfd;
      17'd48143: data = 8'hfc;
      17'd48144: data = 8'hfe;
      17'd48145: data = 8'hfd;
      17'd48146: data = 8'hfe;
      17'd48147: data = 8'hfe;
      17'd48148: data = 8'h00;
      17'd48149: data = 8'h01;
      17'd48150: data = 8'h01;
      17'd48151: data = 8'h01;
      17'd48152: data = 8'h00;
      17'd48153: data = 8'h00;
      17'd48154: data = 8'h00;
      17'd48155: data = 8'hfe;
      17'd48156: data = 8'hfe;
      17'd48157: data = 8'hfd;
      17'd48158: data = 8'hfd;
      17'd48159: data = 8'hfe;
      17'd48160: data = 8'hfe;
      17'd48161: data = 8'hfe;
      17'd48162: data = 8'h01;
      17'd48163: data = 8'h01;
      17'd48164: data = 8'h01;
      17'd48165: data = 8'h02;
      17'd48166: data = 8'h02;
      17'd48167: data = 8'h02;
      17'd48168: data = 8'h00;
      17'd48169: data = 8'hfe;
      17'd48170: data = 8'hfd;
      17'd48171: data = 8'hfd;
      17'd48172: data = 8'hfd;
      17'd48173: data = 8'hfd;
      17'd48174: data = 8'hfd;
      17'd48175: data = 8'hfd;
      17'd48176: data = 8'hfd;
      17'd48177: data = 8'h00;
      17'd48178: data = 8'h01;
      17'd48179: data = 8'h01;
      17'd48180: data = 8'h01;
      17'd48181: data = 8'h01;
      17'd48182: data = 8'h00;
      17'd48183: data = 8'h00;
      17'd48184: data = 8'hfd;
      17'd48185: data = 8'hfd;
      17'd48186: data = 8'hfd;
      17'd48187: data = 8'hfc;
      17'd48188: data = 8'hfc;
      17'd48189: data = 8'hfc;
      17'd48190: data = 8'hfd;
      17'd48191: data = 8'h01;
      17'd48192: data = 8'h00;
      17'd48193: data = 8'h01;
      17'd48194: data = 8'h01;
      17'd48195: data = 8'h00;
      17'd48196: data = 8'h00;
      17'd48197: data = 8'hfe;
      17'd48198: data = 8'h00;
      17'd48199: data = 8'h00;
      17'd48200: data = 8'hfd;
      17'd48201: data = 8'hfd;
      17'd48202: data = 8'hfd;
      17'd48203: data = 8'hfd;
      17'd48204: data = 8'hfe;
      17'd48205: data = 8'hfe;
      17'd48206: data = 8'h00;
      17'd48207: data = 8'h00;
      17'd48208: data = 8'h01;
      17'd48209: data = 8'h01;
      17'd48210: data = 8'h00;
      17'd48211: data = 8'h00;
      17'd48212: data = 8'h00;
      17'd48213: data = 8'h01;
      17'd48214: data = 8'h00;
      17'd48215: data = 8'h01;
      17'd48216: data = 8'h00;
      17'd48217: data = 8'hfe;
      17'd48218: data = 8'hfe;
      17'd48219: data = 8'hfe;
      17'd48220: data = 8'h00;
      17'd48221: data = 8'h01;
      17'd48222: data = 8'h02;
      17'd48223: data = 8'h01;
      17'd48224: data = 8'h01;
      17'd48225: data = 8'h02;
      17'd48226: data = 8'h01;
      17'd48227: data = 8'h00;
      17'd48228: data = 8'h00;
      17'd48229: data = 8'h00;
      17'd48230: data = 8'h00;
      17'd48231: data = 8'h00;
      17'd48232: data = 8'hfe;
      17'd48233: data = 8'hfe;
      17'd48234: data = 8'h00;
      17'd48235: data = 8'h01;
      17'd48236: data = 8'h01;
      17'd48237: data = 8'h02;
      17'd48238: data = 8'h01;
      17'd48239: data = 8'h01;
      17'd48240: data = 8'h01;
      17'd48241: data = 8'hfe;
      17'd48242: data = 8'hfe;
      17'd48243: data = 8'h00;
      17'd48244: data = 8'h00;
      17'd48245: data = 8'hfe;
      17'd48246: data = 8'hfe;
      17'd48247: data = 8'hfe;
      17'd48248: data = 8'hfe;
      17'd48249: data = 8'h00;
      17'd48250: data = 8'h01;
      17'd48251: data = 8'h00;
      17'd48252: data = 8'h01;
      17'd48253: data = 8'h01;
      17'd48254: data = 8'h00;
      17'd48255: data = 8'h00;
      17'd48256: data = 8'hfe;
      17'd48257: data = 8'hfe;
      17'd48258: data = 8'hfe;
      17'd48259: data = 8'hfd;
      17'd48260: data = 8'hfd;
      17'd48261: data = 8'hfd;
      17'd48262: data = 8'hfe;
      17'd48263: data = 8'hfe;
      17'd48264: data = 8'h00;
      17'd48265: data = 8'h00;
      17'd48266: data = 8'h00;
      17'd48267: data = 8'h00;
      17'd48268: data = 8'hfe;
      17'd48269: data = 8'hfe;
      17'd48270: data = 8'hfe;
      17'd48271: data = 8'hfd;
      17'd48272: data = 8'hfd;
      17'd48273: data = 8'hfd;
      17'd48274: data = 8'hfe;
      17'd48275: data = 8'hfe;
      17'd48276: data = 8'h00;
      17'd48277: data = 8'h00;
      17'd48278: data = 8'h00;
      17'd48279: data = 8'h01;
      17'd48280: data = 8'h01;
      17'd48281: data = 8'h00;
      17'd48282: data = 8'h00;
      17'd48283: data = 8'hfe;
      17'd48284: data = 8'hfe;
      17'd48285: data = 8'hfd;
      17'd48286: data = 8'hfc;
      17'd48287: data = 8'hfc;
      17'd48288: data = 8'hfd;
      17'd48289: data = 8'hfe;
      17'd48290: data = 8'hfd;
      17'd48291: data = 8'hfe;
      17'd48292: data = 8'h00;
      17'd48293: data = 8'h00;
      17'd48294: data = 8'h00;
      17'd48295: data = 8'h00;
      17'd48296: data = 8'h00;
      17'd48297: data = 8'h00;
      17'd48298: data = 8'h00;
      17'd48299: data = 8'h00;
      17'd48300: data = 8'hfd;
      17'd48301: data = 8'hfd;
      17'd48302: data = 8'hfd;
      17'd48303: data = 8'hfe;
      17'd48304: data = 8'hfe;
      17'd48305: data = 8'hfe;
      17'd48306: data = 8'hfd;
      17'd48307: data = 8'hfe;
      17'd48308: data = 8'h00;
      17'd48309: data = 8'h01;
      17'd48310: data = 8'h00;
      17'd48311: data = 8'hfe;
      17'd48312: data = 8'hfe;
      17'd48313: data = 8'hfe;
      17'd48314: data = 8'hfd;
      17'd48315: data = 8'hfc;
      17'd48316: data = 8'hfc;
      17'd48317: data = 8'hfd;
      17'd48318: data = 8'hfe;
      17'd48319: data = 8'h00;
      17'd48320: data = 8'h01;
      17'd48321: data = 8'h00;
      17'd48322: data = 8'h01;
      17'd48323: data = 8'h02;
      17'd48324: data = 8'h02;
      17'd48325: data = 8'h00;
      17'd48326: data = 8'h00;
      17'd48327: data = 8'h00;
      17'd48328: data = 8'hfd;
      17'd48329: data = 8'hfd;
      17'd48330: data = 8'hfd;
      17'd48331: data = 8'hfd;
      17'd48332: data = 8'hfd;
      17'd48333: data = 8'hfd;
      17'd48334: data = 8'hfe;
      17'd48335: data = 8'h00;
      17'd48336: data = 8'h01;
      17'd48337: data = 8'h02;
      17'd48338: data = 8'h01;
      17'd48339: data = 8'h01;
      17'd48340: data = 8'h01;
      17'd48341: data = 8'h00;
      17'd48342: data = 8'h00;
      17'd48343: data = 8'h00;
      17'd48344: data = 8'hfe;
      17'd48345: data = 8'hfe;
      17'd48346: data = 8'h00;
      17'd48347: data = 8'h00;
      17'd48348: data = 8'h00;
      17'd48349: data = 8'h00;
      17'd48350: data = 8'hfe;
      17'd48351: data = 8'h01;
      17'd48352: data = 8'h01;
      17'd48353: data = 8'h01;
      17'd48354: data = 8'h00;
      17'd48355: data = 8'hfe;
      17'd48356: data = 8'h01;
      17'd48357: data = 8'hfe;
      17'd48358: data = 8'hfe;
      17'd48359: data = 8'hfd;
      17'd48360: data = 8'hfc;
      17'd48361: data = 8'hfe;
      17'd48362: data = 8'hfe;
      17'd48363: data = 8'hfe;
      17'd48364: data = 8'h00;
      17'd48365: data = 8'h00;
      17'd48366: data = 8'h01;
      17'd48367: data = 8'h01;
      17'd48368: data = 8'h00;
      17'd48369: data = 8'h00;
      17'd48370: data = 8'hfe;
      17'd48371: data = 8'h00;
      17'd48372: data = 8'hfe;
      17'd48373: data = 8'hfd;
      17'd48374: data = 8'hfe;
      17'd48375: data = 8'hfe;
      17'd48376: data = 8'h00;
      17'd48377: data = 8'hfe;
      17'd48378: data = 8'h00;
      17'd48379: data = 8'h00;
      17'd48380: data = 8'h01;
      17'd48381: data = 8'h01;
      17'd48382: data = 8'h00;
      17'd48383: data = 8'hfe;
      17'd48384: data = 8'hfe;
      17'd48385: data = 8'h00;
      17'd48386: data = 8'hfd;
      17'd48387: data = 8'hfd;
      17'd48388: data = 8'hfd;
      17'd48389: data = 8'hfe;
      17'd48390: data = 8'hfd;
      17'd48391: data = 8'hfe;
      17'd48392: data = 8'h01;
      17'd48393: data = 8'h00;
      17'd48394: data = 8'h01;
      17'd48395: data = 8'h02;
      17'd48396: data = 8'h01;
      17'd48397: data = 8'h02;
      17'd48398: data = 8'h01;
      17'd48399: data = 8'h01;
      17'd48400: data = 8'h00;
      17'd48401: data = 8'h00;
      17'd48402: data = 8'hfe;
      17'd48403: data = 8'hfd;
      17'd48404: data = 8'h00;
      17'd48405: data = 8'hfd;
      17'd48406: data = 8'h00;
      17'd48407: data = 8'h00;
      17'd48408: data = 8'h00;
      17'd48409: data = 8'h02;
      17'd48410: data = 8'h01;
      17'd48411: data = 8'h01;
      17'd48412: data = 8'h02;
      17'd48413: data = 8'h01;
      17'd48414: data = 8'h00;
      17'd48415: data = 8'h00;
      17'd48416: data = 8'hfe;
      17'd48417: data = 8'hfd;
      17'd48418: data = 8'hfd;
      17'd48419: data = 8'hfd;
      17'd48420: data = 8'hfe;
      17'd48421: data = 8'hfe;
      17'd48422: data = 8'h01;
      17'd48423: data = 8'h01;
      17'd48424: data = 8'h01;
      17'd48425: data = 8'h01;
      17'd48426: data = 8'h01;
      17'd48427: data = 8'h01;
      17'd48428: data = 8'h00;
      17'd48429: data = 8'h00;
      17'd48430: data = 8'hfe;
      17'd48431: data = 8'hfe;
      17'd48432: data = 8'hfe;
      17'd48433: data = 8'hfe;
      17'd48434: data = 8'hfd;
      17'd48435: data = 8'hfd;
      17'd48436: data = 8'h00;
      17'd48437: data = 8'hfe;
      17'd48438: data = 8'h00;
      17'd48439: data = 8'h00;
      17'd48440: data = 8'h00;
      17'd48441: data = 8'h00;
      17'd48442: data = 8'h00;
      17'd48443: data = 8'hfe;
      17'd48444: data = 8'hfe;
      17'd48445: data = 8'hfe;
      17'd48446: data = 8'hfd;
      17'd48447: data = 8'hfd;
      17'd48448: data = 8'hfd;
      17'd48449: data = 8'hfd;
      17'd48450: data = 8'hfd;
      17'd48451: data = 8'hfe;
      17'd48452: data = 8'hfe;
      17'd48453: data = 8'h00;
      17'd48454: data = 8'h00;
      17'd48455: data = 8'h00;
      17'd48456: data = 8'h00;
      17'd48457: data = 8'h00;
      17'd48458: data = 8'h01;
      17'd48459: data = 8'h00;
      17'd48460: data = 8'h00;
      17'd48461: data = 8'hfe;
      17'd48462: data = 8'hfe;
      17'd48463: data = 8'h00;
      17'd48464: data = 8'h00;
      17'd48465: data = 8'h00;
      17'd48466: data = 8'h00;
      17'd48467: data = 8'h00;
      17'd48468: data = 8'h00;
      17'd48469: data = 8'h00;
      17'd48470: data = 8'h01;
      17'd48471: data = 8'h01;
      17'd48472: data = 8'h00;
      17'd48473: data = 8'h00;
      17'd48474: data = 8'hfe;
      17'd48475: data = 8'hfe;
      17'd48476: data = 8'hfe;
      17'd48477: data = 8'hfe;
      17'd48478: data = 8'hfe;
      17'd48479: data = 8'hfe;
      17'd48480: data = 8'hfe;
      17'd48481: data = 8'hfe;
      17'd48482: data = 8'h00;
      17'd48483: data = 8'h01;
      17'd48484: data = 8'h01;
      17'd48485: data = 8'hfe;
      17'd48486: data = 8'hfe;
      17'd48487: data = 8'h00;
      17'd48488: data = 8'h01;
      17'd48489: data = 8'h00;
      17'd48490: data = 8'hfe;
      17'd48491: data = 8'h00;
      17'd48492: data = 8'h00;
      17'd48493: data = 8'hfe;
      17'd48494: data = 8'h00;
      17'd48495: data = 8'h00;
      17'd48496: data = 8'hfe;
      17'd48497: data = 8'hfe;
      17'd48498: data = 8'hfe;
      17'd48499: data = 8'h00;
      17'd48500: data = 8'h00;
      17'd48501: data = 8'h00;
      17'd48502: data = 8'h01;
      17'd48503: data = 8'h01;
      17'd48504: data = 8'h00;
      17'd48505: data = 8'h00;
      17'd48506: data = 8'h00;
      17'd48507: data = 8'hfe;
      17'd48508: data = 8'hfe;
      17'd48509: data = 8'hfe;
      17'd48510: data = 8'h00;
      17'd48511: data = 8'h00;
      17'd48512: data = 8'hfd;
      17'd48513: data = 8'hfe;
      17'd48514: data = 8'h00;
      17'd48515: data = 8'h01;
      17'd48516: data = 8'h01;
      17'd48517: data = 8'hfe;
      17'd48518: data = 8'h00;
      17'd48519: data = 8'h01;
      17'd48520: data = 8'h00;
      17'd48521: data = 8'hfe;
      17'd48522: data = 8'hfe;
      17'd48523: data = 8'hfe;
      17'd48524: data = 8'h00;
      17'd48525: data = 8'h00;
      17'd48526: data = 8'hfe;
      17'd48527: data = 8'h00;
      17'd48528: data = 8'h00;
      17'd48529: data = 8'h00;
      17'd48530: data = 8'h00;
      17'd48531: data = 8'h00;
      17'd48532: data = 8'h01;
      17'd48533: data = 8'h01;
      17'd48534: data = 8'h01;
      17'd48535: data = 8'h00;
      17'd48536: data = 8'h00;
      17'd48537: data = 8'h00;
      17'd48538: data = 8'h00;
      17'd48539: data = 8'hfe;
      17'd48540: data = 8'h00;
      17'd48541: data = 8'hfe;
      17'd48542: data = 8'hfe;
      17'd48543: data = 8'hfe;
      17'd48544: data = 8'h00;
      17'd48545: data = 8'h00;
      17'd48546: data = 8'h00;
      17'd48547: data = 8'h01;
      17'd48548: data = 8'h00;
      17'd48549: data = 8'h01;
      17'd48550: data = 8'h01;
      17'd48551: data = 8'h01;
      17'd48552: data = 8'hfe;
      17'd48553: data = 8'hfe;
      17'd48554: data = 8'h00;
      17'd48555: data = 8'h00;
      17'd48556: data = 8'h02;
      17'd48557: data = 8'h00;
      17'd48558: data = 8'hfe;
      17'd48559: data = 8'h00;
      17'd48560: data = 8'h01;
      17'd48561: data = 8'h01;
      17'd48562: data = 8'h00;
      17'd48563: data = 8'h00;
      17'd48564: data = 8'h01;
      17'd48565: data = 8'h02;
      17'd48566: data = 8'h01;
      17'd48567: data = 8'h01;
      17'd48568: data = 8'h01;
      17'd48569: data = 8'h01;
      17'd48570: data = 8'h01;
      17'd48571: data = 8'h01;
      17'd48572: data = 8'h00;
      17'd48573: data = 8'h00;
      17'd48574: data = 8'h00;
      17'd48575: data = 8'h00;
      17'd48576: data = 8'h00;
      17'd48577: data = 8'h00;
      17'd48578: data = 8'h01;
      17'd48579: data = 8'h01;
      17'd48580: data = 8'h01;
      17'd48581: data = 8'h01;
      17'd48582: data = 8'h01;
      17'd48583: data = 8'h01;
      17'd48584: data = 8'h00;
      17'd48585: data = 8'h00;
      17'd48586: data = 8'h01;
      17'd48587: data = 8'h01;
      17'd48588: data = 8'h00;
      17'd48589: data = 8'h00;
      17'd48590: data = 8'hfe;
      17'd48591: data = 8'h00;
      17'd48592: data = 8'h00;
      17'd48593: data = 8'h00;
      17'd48594: data = 8'h00;
      17'd48595: data = 8'h01;
      17'd48596: data = 8'h01;
      17'd48597: data = 8'h01;
      17'd48598: data = 8'h01;
      17'd48599: data = 8'h00;
      17'd48600: data = 8'h01;
      17'd48601: data = 8'h00;
      17'd48602: data = 8'hfe;
      17'd48603: data = 8'hfe;
      17'd48604: data = 8'hfe;
      17'd48605: data = 8'hfe;
      17'd48606: data = 8'hfe;
      17'd48607: data = 8'hfd;
      17'd48608: data = 8'hfd;
      17'd48609: data = 8'h00;
      17'd48610: data = 8'h01;
      17'd48611: data = 8'h00;
      17'd48612: data = 8'h00;
      17'd48613: data = 8'h00;
      17'd48614: data = 8'h00;
      17'd48615: data = 8'h00;
      17'd48616: data = 8'h00;
      17'd48617: data = 8'hfe;
      17'd48618: data = 8'hfe;
      17'd48619: data = 8'hfe;
      17'd48620: data = 8'hfd;
      17'd48621: data = 8'hfd;
      17'd48622: data = 8'hfc;
      17'd48623: data = 8'hfe;
      17'd48624: data = 8'hfe;
      17'd48625: data = 8'hfe;
      17'd48626: data = 8'hfe;
      17'd48627: data = 8'h00;
      17'd48628: data = 8'h00;
      17'd48629: data = 8'h01;
      17'd48630: data = 8'h01;
      17'd48631: data = 8'h01;
      17'd48632: data = 8'h00;
      17'd48633: data = 8'h00;
      17'd48634: data = 8'h00;
      17'd48635: data = 8'hfd;
      17'd48636: data = 8'hfd;
      17'd48637: data = 8'hfd;
      17'd48638: data = 8'hfe;
      17'd48639: data = 8'hfe;
      17'd48640: data = 8'hfe;
      17'd48641: data = 8'hfe;
      17'd48642: data = 8'h00;
      17'd48643: data = 8'h00;
      17'd48644: data = 8'h00;
      17'd48645: data = 8'h00;
      17'd48646: data = 8'h00;
      17'd48647: data = 8'h01;
      17'd48648: data = 8'hfe;
      17'd48649: data = 8'hfe;
      17'd48650: data = 8'h00;
      17'd48651: data = 8'hfe;
      17'd48652: data = 8'hfd;
      17'd48653: data = 8'hfd;
      17'd48654: data = 8'hfe;
      17'd48655: data = 8'hfe;
      17'd48656: data = 8'hfe;
      17'd48657: data = 8'h00;
      17'd48658: data = 8'hfe;
      17'd48659: data = 8'h00;
      17'd48660: data = 8'h01;
      17'd48661: data = 8'h01;
      17'd48662: data = 8'h02;
      17'd48663: data = 8'h01;
      17'd48664: data = 8'hfe;
      17'd48665: data = 8'hfe;
      17'd48666: data = 8'h00;
      17'd48667: data = 8'hfe;
      17'd48668: data = 8'hfe;
      17'd48669: data = 8'hfe;
      17'd48670: data = 8'hfe;
      17'd48671: data = 8'hfe;
      17'd48672: data = 8'hfe;
      17'd48673: data = 8'hfe;
      17'd48674: data = 8'h00;
      17'd48675: data = 8'h00;
      17'd48676: data = 8'hfe;
      17'd48677: data = 8'h00;
      17'd48678: data = 8'h01;
      17'd48679: data = 8'h01;
      17'd48680: data = 8'h00;
      17'd48681: data = 8'h00;
      17'd48682: data = 8'h00;
      17'd48683: data = 8'hfe;
      17'd48684: data = 8'h00;
      17'd48685: data = 8'hfd;
      17'd48686: data = 8'hfe;
      17'd48687: data = 8'hfd;
      17'd48688: data = 8'hfd;
      17'd48689: data = 8'hfe;
      17'd48690: data = 8'hfe;
      17'd48691: data = 8'h01;
      17'd48692: data = 8'hfe;
      17'd48693: data = 8'h01;
      17'd48694: data = 8'h02;
      17'd48695: data = 8'h01;
      17'd48696: data = 8'h01;
      17'd48697: data = 8'hfe;
      17'd48698: data = 8'h00;
      17'd48699: data = 8'hfe;
      17'd48700: data = 8'hfe;
      17'd48701: data = 8'hfe;
      17'd48702: data = 8'hfd;
      17'd48703: data = 8'hfe;
      17'd48704: data = 8'h00;
      17'd48705: data = 8'hfe;
      17'd48706: data = 8'hfe;
      17'd48707: data = 8'hfe;
      17'd48708: data = 8'h00;
      17'd48709: data = 8'h00;
      17'd48710: data = 8'h01;
      17'd48711: data = 8'h00;
      17'd48712: data = 8'h00;
      17'd48713: data = 8'hfe;
      17'd48714: data = 8'hfd;
      17'd48715: data = 8'hfd;
      17'd48716: data = 8'hfe;
      17'd48717: data = 8'hfe;
      17'd48718: data = 8'hfd;
      17'd48719: data = 8'hfd;
      17'd48720: data = 8'h00;
      17'd48721: data = 8'h00;
      17'd48722: data = 8'hfe;
      17'd48723: data = 8'h01;
      17'd48724: data = 8'h01;
      17'd48725: data = 8'h01;
      17'd48726: data = 8'h01;
      17'd48727: data = 8'h01;
      17'd48728: data = 8'h01;
      17'd48729: data = 8'hfe;
      17'd48730: data = 8'hfd;
      17'd48731: data = 8'hfe;
      17'd48732: data = 8'hfe;
      17'd48733: data = 8'hfd;
      17'd48734: data = 8'hfe;
      17'd48735: data = 8'hfd;
      17'd48736: data = 8'hfe;
      17'd48737: data = 8'hfe;
      17'd48738: data = 8'hfe;
      17'd48739: data = 8'hfe;
      17'd48740: data = 8'h00;
      17'd48741: data = 8'h01;
      17'd48742: data = 8'h00;
      17'd48743: data = 8'h00;
      17'd48744: data = 8'hfe;
      17'd48745: data = 8'hfd;
      17'd48746: data = 8'hfd;
      17'd48747: data = 8'hfe;
      17'd48748: data = 8'hfc;
      17'd48749: data = 8'hfa;
      17'd48750: data = 8'hfc;
      17'd48751: data = 8'hfe;
      17'd48752: data = 8'hfe;
      17'd48753: data = 8'hfd;
      17'd48754: data = 8'h00;
      17'd48755: data = 8'hfe;
      17'd48756: data = 8'h00;
      17'd48757: data = 8'h00;
      17'd48758: data = 8'hfe;
      17'd48759: data = 8'h00;
      17'd48760: data = 8'hfe;
      17'd48761: data = 8'hfe;
      17'd48762: data = 8'hfd;
      17'd48763: data = 8'hfd;
      17'd48764: data = 8'hfd;
      17'd48765: data = 8'hfc;
      17'd48766: data = 8'hfd;
      17'd48767: data = 8'hfd;
      17'd48768: data = 8'hfe;
      17'd48769: data = 8'h00;
      17'd48770: data = 8'h00;
      17'd48771: data = 8'h00;
      17'd48772: data = 8'h01;
      17'd48773: data = 8'h01;
      17'd48774: data = 8'hfe;
      17'd48775: data = 8'hfe;
      17'd48776: data = 8'hfe;
      17'd48777: data = 8'hfc;
      17'd48778: data = 8'hfc;
      17'd48779: data = 8'hfd;
      17'd48780: data = 8'hfd;
      17'd48781: data = 8'hfd;
      17'd48782: data = 8'hfe;
      17'd48783: data = 8'hfe;
      17'd48784: data = 8'h00;
      17'd48785: data = 8'hfe;
      17'd48786: data = 8'hfe;
      17'd48787: data = 8'hfe;
      17'd48788: data = 8'h00;
      17'd48789: data = 8'h01;
      17'd48790: data = 8'h00;
      17'd48791: data = 8'hfe;
      17'd48792: data = 8'h00;
      17'd48793: data = 8'h00;
      17'd48794: data = 8'hfe;
      17'd48795: data = 8'hfe;
      17'd48796: data = 8'hfe;
      17'd48797: data = 8'hfe;
      17'd48798: data = 8'hfe;
      17'd48799: data = 8'hfe;
      17'd48800: data = 8'hfe;
      17'd48801: data = 8'hfe;
      17'd48802: data = 8'hfe;
      17'd48803: data = 8'hfe;
      17'd48804: data = 8'hfe;
      17'd48805: data = 8'hfe;
      17'd48806: data = 8'h00;
      17'd48807: data = 8'hfe;
      17'd48808: data = 8'hfe;
      17'd48809: data = 8'h00;
      17'd48810: data = 8'h00;
      17'd48811: data = 8'h00;
      17'd48812: data = 8'h00;
      17'd48813: data = 8'hfe;
      17'd48814: data = 8'hfe;
      17'd48815: data = 8'hfe;
      17'd48816: data = 8'h00;
      17'd48817: data = 8'hfe;
      17'd48818: data = 8'h00;
      17'd48819: data = 8'h00;
      17'd48820: data = 8'hfe;
      17'd48821: data = 8'h00;
      17'd48822: data = 8'hfe;
      17'd48823: data = 8'h00;
      17'd48824: data = 8'h00;
      17'd48825: data = 8'h01;
      17'd48826: data = 8'h01;
      17'd48827: data = 8'h01;
      17'd48828: data = 8'h01;
      17'd48829: data = 8'h01;
      17'd48830: data = 8'h01;
      17'd48831: data = 8'h00;
      17'd48832: data = 8'h00;
      17'd48833: data = 8'hfe;
      17'd48834: data = 8'h00;
      17'd48835: data = 8'h00;
      17'd48836: data = 8'h02;
      17'd48837: data = 8'h01;
      17'd48838: data = 8'h00;
      17'd48839: data = 8'h02;
      17'd48840: data = 8'h02;
      17'd48841: data = 8'h01;
      17'd48842: data = 8'h01;
      17'd48843: data = 8'h00;
      17'd48844: data = 8'hfe;
      17'd48845: data = 8'hfe;
      17'd48846: data = 8'hfd;
      17'd48847: data = 8'hfe;
      17'd48848: data = 8'hfe;
      17'd48849: data = 8'hfd;
      17'd48850: data = 8'hfe;
      17'd48851: data = 8'h00;
      17'd48852: data = 8'hfe;
      17'd48853: data = 8'h00;
      17'd48854: data = 8'h01;
      17'd48855: data = 8'h01;
      17'd48856: data = 8'h02;
      17'd48857: data = 8'h01;
      17'd48858: data = 8'h01;
      17'd48859: data = 8'h00;
      17'd48860: data = 8'h00;
      17'd48861: data = 8'h00;
      17'd48862: data = 8'hfd;
      17'd48863: data = 8'hfe;
      17'd48864: data = 8'hfe;
      17'd48865: data = 8'hfd;
      17'd48866: data = 8'h00;
      17'd48867: data = 8'h00;
      17'd48868: data = 8'h01;
      17'd48869: data = 8'h00;
      17'd48870: data = 8'h00;
      17'd48871: data = 8'h01;
      17'd48872: data = 8'h01;
      17'd48873: data = 8'h01;
      17'd48874: data = 8'hfe;
      17'd48875: data = 8'hfe;
      17'd48876: data = 8'hfe;
      17'd48877: data = 8'hfd;
      17'd48878: data = 8'hfd;
      17'd48879: data = 8'hfd;
      17'd48880: data = 8'hfe;
      17'd48881: data = 8'hfe;
      17'd48882: data = 8'h00;
      17'd48883: data = 8'h01;
      17'd48884: data = 8'h02;
      17'd48885: data = 8'h01;
      17'd48886: data = 8'h01;
      17'd48887: data = 8'h02;
      17'd48888: data = 8'h01;
      17'd48889: data = 8'h01;
      17'd48890: data = 8'h01;
      17'd48891: data = 8'h00;
      17'd48892: data = 8'hfe;
      17'd48893: data = 8'hfd;
      17'd48894: data = 8'hfe;
      17'd48895: data = 8'hfe;
      17'd48896: data = 8'hfe;
      17'd48897: data = 8'h00;
      17'd48898: data = 8'h01;
      17'd48899: data = 8'h01;
      17'd48900: data = 8'h00;
      17'd48901: data = 8'h02;
      17'd48902: data = 8'h02;
      17'd48903: data = 8'h00;
      17'd48904: data = 8'h01;
      17'd48905: data = 8'h00;
      17'd48906: data = 8'hfe;
      17'd48907: data = 8'hfe;
      17'd48908: data = 8'hfd;
      17'd48909: data = 8'hfe;
      17'd48910: data = 8'hfe;
      17'd48911: data = 8'hfe;
      17'd48912: data = 8'h00;
      17'd48913: data = 8'h00;
      17'd48914: data = 8'h00;
      17'd48915: data = 8'h01;
      17'd48916: data = 8'h01;
      17'd48917: data = 8'h01;
      17'd48918: data = 8'h01;
      17'd48919: data = 8'h00;
      17'd48920: data = 8'h00;
      17'd48921: data = 8'h00;
      17'd48922: data = 8'hfd;
      17'd48923: data = 8'hfe;
      17'd48924: data = 8'hfe;
      17'd48925: data = 8'hfe;
      17'd48926: data = 8'h00;
      17'd48927: data = 8'h02;
      17'd48928: data = 8'h00;
      17'd48929: data = 8'h01;
      17'd48930: data = 8'h00;
      17'd48931: data = 8'h00;
      17'd48932: data = 8'h01;
      17'd48933: data = 8'hfe;
      17'd48934: data = 8'hfe;
      17'd48935: data = 8'hfe;
      17'd48936: data = 8'hfe;
      17'd48937: data = 8'hfe;
      17'd48938: data = 8'hfe;
      17'd48939: data = 8'h00;
      17'd48940: data = 8'hfe;
      17'd48941: data = 8'h00;
      17'd48942: data = 8'h00;
      17'd48943: data = 8'h00;
      17'd48944: data = 8'h00;
      17'd48945: data = 8'h00;
      17'd48946: data = 8'hfe;
      17'd48947: data = 8'hfe;
      17'd48948: data = 8'hfe;
      17'd48949: data = 8'hfd;
      17'd48950: data = 8'hfd;
      17'd48951: data = 8'hfd;
      17'd48952: data = 8'hfe;
      17'd48953: data = 8'hfd;
      17'd48954: data = 8'hfe;
      17'd48955: data = 8'h00;
      17'd48956: data = 8'h00;
      17'd48957: data = 8'h01;
      17'd48958: data = 8'h01;
      17'd48959: data = 8'h01;
      17'd48960: data = 8'h00;
      17'd48961: data = 8'h00;
      17'd48962: data = 8'hfe;
      17'd48963: data = 8'hfd;
      17'd48964: data = 8'hfd;
      17'd48965: data = 8'hfd;
      17'd48966: data = 8'hfd;
      17'd48967: data = 8'hfe;
      17'd48968: data = 8'hfe;
      17'd48969: data = 8'hfe;
      17'd48970: data = 8'h00;
      17'd48971: data = 8'h00;
      17'd48972: data = 8'h01;
      17'd48973: data = 8'h00;
      17'd48974: data = 8'h00;
      17'd48975: data = 8'hfe;
      17'd48976: data = 8'hfe;
      17'd48977: data = 8'hfe;
      17'd48978: data = 8'hfd;
      17'd48979: data = 8'hfd;
      17'd48980: data = 8'hfc;
      17'd48981: data = 8'hfd;
      17'd48982: data = 8'hfd;
      17'd48983: data = 8'hfe;
      17'd48984: data = 8'h00;
      17'd48985: data = 8'h00;
      17'd48986: data = 8'h00;
      17'd48987: data = 8'h01;
      17'd48988: data = 8'h00;
      17'd48989: data = 8'hfe;
      17'd48990: data = 8'hfe;
      17'd48991: data = 8'hfe;
      17'd48992: data = 8'hfc;
      17'd48993: data = 8'hfc;
      17'd48994: data = 8'hfd;
      17'd48995: data = 8'hfc;
      17'd48996: data = 8'hfc;
      17'd48997: data = 8'hfd;
      17'd48998: data = 8'hfe;
      17'd48999: data = 8'h00;
      17'd49000: data = 8'h01;
      17'd49001: data = 8'h01;
      17'd49002: data = 8'h01;
      17'd49003: data = 8'h00;
      17'd49004: data = 8'h00;
      17'd49005: data = 8'h00;
      17'd49006: data = 8'hfd;
      17'd49007: data = 8'hfa;
      17'd49008: data = 8'hfd;
      17'd49009: data = 8'hfd;
      17'd49010: data = 8'hfd;
      17'd49011: data = 8'hfe;
      17'd49012: data = 8'h00;
      17'd49013: data = 8'h01;
      17'd49014: data = 8'h00;
      17'd49015: data = 8'h01;
      17'd49016: data = 8'h01;
      17'd49017: data = 8'h00;
      17'd49018: data = 8'h00;
      17'd49019: data = 8'hfe;
      17'd49020: data = 8'hfd;
      17'd49021: data = 8'hfd;
      17'd49022: data = 8'hfd;
      17'd49023: data = 8'hfc;
      17'd49024: data = 8'hfd;
      17'd49025: data = 8'hfe;
      17'd49026: data = 8'hfe;
      17'd49027: data = 8'hfe;
      17'd49028: data = 8'h00;
      17'd49029: data = 8'h01;
      17'd49030: data = 8'h01;
      17'd49031: data = 8'h02;
      17'd49032: data = 8'h01;
      17'd49033: data = 8'hfe;
      17'd49034: data = 8'hfe;
      17'd49035: data = 8'hfe;
      17'd49036: data = 8'hfc;
      17'd49037: data = 8'hfc;
      17'd49038: data = 8'hfd;
      17'd49039: data = 8'hfc;
      17'd49040: data = 8'hfe;
      17'd49041: data = 8'hfd;
      17'd49042: data = 8'hfe;
      17'd49043: data = 8'h00;
      17'd49044: data = 8'h00;
      17'd49045: data = 8'h00;
      17'd49046: data = 8'h00;
      17'd49047: data = 8'hfe;
      17'd49048: data = 8'hfe;
      17'd49049: data = 8'hfe;
      17'd49050: data = 8'hfd;
      17'd49051: data = 8'hfe;
      17'd49052: data = 8'hfd;
      17'd49053: data = 8'hfd;
      17'd49054: data = 8'hfc;
      17'd49055: data = 8'hfe;
      17'd49056: data = 8'hfe;
      17'd49057: data = 8'hfe;
      17'd49058: data = 8'h01;
      17'd49059: data = 8'h00;
      17'd49060: data = 8'h00;
      17'd49061: data = 8'h01;
      17'd49062: data = 8'h00;
      17'd49063: data = 8'h00;
      17'd49064: data = 8'h00;
      17'd49065: data = 8'hfd;
      17'd49066: data = 8'hfd;
      17'd49067: data = 8'hfe;
      17'd49068: data = 8'hfd;
      17'd49069: data = 8'h01;
      17'd49070: data = 8'h00;
      17'd49071: data = 8'hfe;
      17'd49072: data = 8'h00;
      17'd49073: data = 8'h01;
      17'd49074: data = 8'h01;
      17'd49075: data = 8'h01;
      17'd49076: data = 8'h00;
      17'd49077: data = 8'h00;
      17'd49078: data = 8'h00;
      17'd49079: data = 8'hfe;
      17'd49080: data = 8'hfe;
      17'd49081: data = 8'hfe;
      17'd49082: data = 8'hfe;
      17'd49083: data = 8'hfe;
      17'd49084: data = 8'hfe;
      17'd49085: data = 8'h01;
      17'd49086: data = 8'h01;
      17'd49087: data = 8'h01;
      17'd49088: data = 8'h01;
      17'd49089: data = 8'h02;
      17'd49090: data = 8'h01;
      17'd49091: data = 8'h00;
      17'd49092: data = 8'h00;
      17'd49093: data = 8'hfe;
      17'd49094: data = 8'h00;
      17'd49095: data = 8'hfe;
      17'd49096: data = 8'hfd;
      17'd49097: data = 8'h00;
      17'd49098: data = 8'h01;
      17'd49099: data = 8'h00;
      17'd49100: data = 8'h00;
      17'd49101: data = 8'h00;
      17'd49102: data = 8'hfe;
      17'd49103: data = 8'h00;
      17'd49104: data = 8'h00;
      17'd49105: data = 8'h00;
      17'd49106: data = 8'h00;
      17'd49107: data = 8'hfe;
      17'd49108: data = 8'h00;
      17'd49109: data = 8'hfe;
      17'd49110: data = 8'hfe;
      17'd49111: data = 8'h00;
      17'd49112: data = 8'h00;
      17'd49113: data = 8'h00;
      17'd49114: data = 8'h01;
      17'd49115: data = 8'h01;
      17'd49116: data = 8'h00;
      17'd49117: data = 8'h00;
      17'd49118: data = 8'hfe;
      17'd49119: data = 8'hfe;
      17'd49120: data = 8'h00;
      17'd49121: data = 8'h00;
      17'd49122: data = 8'hfe;
      17'd49123: data = 8'h00;
      17'd49124: data = 8'h00;
      17'd49125: data = 8'h00;
      17'd49126: data = 8'h00;
      17'd49127: data = 8'h00;
      17'd49128: data = 8'h00;
      17'd49129: data = 8'hfe;
      17'd49130: data = 8'h00;
      17'd49131: data = 8'h00;
      17'd49132: data = 8'hfe;
      17'd49133: data = 8'hfe;
      17'd49134: data = 8'hfe;
      17'd49135: data = 8'h00;
      17'd49136: data = 8'h00;
      17'd49137: data = 8'h00;
      17'd49138: data = 8'h00;
      17'd49139: data = 8'h00;
      17'd49140: data = 8'h01;
      17'd49141: data = 8'h00;
      17'd49142: data = 8'h00;
      17'd49143: data = 8'h00;
      17'd49144: data = 8'hfe;
      17'd49145: data = 8'hfe;
      17'd49146: data = 8'hfe;
      17'd49147: data = 8'hfd;
      17'd49148: data = 8'hfe;
      17'd49149: data = 8'h00;
      17'd49150: data = 8'hfe;
      17'd49151: data = 8'h01;
      17'd49152: data = 8'h01;
      17'd49153: data = 8'h00;
      17'd49154: data = 8'h01;
      17'd49155: data = 8'h01;
      17'd49156: data = 8'hfe;
      17'd49157: data = 8'hfe;
      17'd49158: data = 8'hfe;
      17'd49159: data = 8'hfc;
      17'd49160: data = 8'hfd;
      17'd49161: data = 8'hfe;
      17'd49162: data = 8'hfd;
      17'd49163: data = 8'hfd;
      17'd49164: data = 8'h01;
      17'd49165: data = 8'h01;
      17'd49166: data = 8'h01;
      17'd49167: data = 8'h02;
      17'd49168: data = 8'h02;
      17'd49169: data = 8'h01;
      17'd49170: data = 8'h00;
      17'd49171: data = 8'h01;
      17'd49172: data = 8'hfe;
      17'd49173: data = 8'hfd;
      17'd49174: data = 8'hfc;
      17'd49175: data = 8'hfc;
      17'd49176: data = 8'hfc;
      17'd49177: data = 8'hfd;
      17'd49178: data = 8'hfe;
      17'd49179: data = 8'hfe;
      17'd49180: data = 8'h00;
      17'd49181: data = 8'h01;
      17'd49182: data = 8'h01;
      17'd49183: data = 8'h01;
      17'd49184: data = 8'h01;
      17'd49185: data = 8'h01;
      17'd49186: data = 8'hfe;
      17'd49187: data = 8'hfe;
      17'd49188: data = 8'hfe;
      17'd49189: data = 8'hfd;
      17'd49190: data = 8'hfd;
      17'd49191: data = 8'hfd;
      17'd49192: data = 8'hfd;
      17'd49193: data = 8'h00;
      17'd49194: data = 8'h01;
      17'd49195: data = 8'h02;
      17'd49196: data = 8'h02;
      17'd49197: data = 8'h04;
      17'd49198: data = 8'h04;
      17'd49199: data = 8'h04;
      17'd49200: data = 8'h02;
      17'd49201: data = 8'hfe;
      17'd49202: data = 8'hfe;
      17'd49203: data = 8'h00;
      17'd49204: data = 8'hfc;
      17'd49205: data = 8'hfc;
      17'd49206: data = 8'hfd;
      17'd49207: data = 8'hfd;
      17'd49208: data = 8'hfe;
      17'd49209: data = 8'h00;
      17'd49210: data = 8'h01;
      17'd49211: data = 8'h02;
      17'd49212: data = 8'h04;
      17'd49213: data = 8'h04;
      17'd49214: data = 8'h02;
      17'd49215: data = 8'h00;
      17'd49216: data = 8'hfe;
      17'd49217: data = 8'hfd;
      17'd49218: data = 8'hfd;
      17'd49219: data = 8'hfe;
      17'd49220: data = 8'hfd;
      17'd49221: data = 8'hfd;
      17'd49222: data = 8'h00;
      17'd49223: data = 8'h00;
      17'd49224: data = 8'h02;
      17'd49225: data = 8'h02;
      17'd49226: data = 8'h02;
      17'd49227: data = 8'h04;
      17'd49228: data = 8'h02;
      17'd49229: data = 8'h02;
      17'd49230: data = 8'h00;
      17'd49231: data = 8'h00;
      17'd49232: data = 8'hfe;
      17'd49233: data = 8'hfe;
      17'd49234: data = 8'hfd;
      17'd49235: data = 8'hfd;
      17'd49236: data = 8'hfe;
      17'd49237: data = 8'hfe;
      17'd49238: data = 8'h01;
      17'd49239: data = 8'h01;
      17'd49240: data = 8'h01;
      17'd49241: data = 8'h01;
      17'd49242: data = 8'h01;
      17'd49243: data = 8'h00;
      17'd49244: data = 8'h00;
      17'd49245: data = 8'h00;
      17'd49246: data = 8'hfe;
      17'd49247: data = 8'hfd;
      17'd49248: data = 8'hfd;
      17'd49249: data = 8'hfe;
      17'd49250: data = 8'hfe;
      17'd49251: data = 8'h00;
      17'd49252: data = 8'h01;
      17'd49253: data = 8'h01;
      17'd49254: data = 8'h04;
      17'd49255: data = 8'h02;
      17'd49256: data = 8'h04;
      17'd49257: data = 8'h01;
      17'd49258: data = 8'h00;
      17'd49259: data = 8'h00;
      17'd49260: data = 8'hfe;
      17'd49261: data = 8'hfe;
      17'd49262: data = 8'hfe;
      17'd49263: data = 8'hfe;
      17'd49264: data = 8'hfe;
      17'd49265: data = 8'hfe;
      17'd49266: data = 8'h00;
      17'd49267: data = 8'h01;
      17'd49268: data = 8'h01;
      17'd49269: data = 8'h01;
      17'd49270: data = 8'h02;
      17'd49271: data = 8'h02;
      17'd49272: data = 8'h00;
      17'd49273: data = 8'h00;
      17'd49274: data = 8'hfe;
      17'd49275: data = 8'hfd;
      17'd49276: data = 8'hfc;
      17'd49277: data = 8'hfc;
      17'd49278: data = 8'hfd;
      17'd49279: data = 8'hfd;
      17'd49280: data = 8'hfd;
      17'd49281: data = 8'h00;
      17'd49282: data = 8'h01;
      17'd49283: data = 8'h01;
      17'd49284: data = 8'h01;
      17'd49285: data = 8'h01;
      17'd49286: data = 8'h01;
      17'd49287: data = 8'h00;
      17'd49288: data = 8'h00;
      17'd49289: data = 8'hfe;
      17'd49290: data = 8'hfd;
      17'd49291: data = 8'hfd;
      17'd49292: data = 8'hfc;
      17'd49293: data = 8'hfc;
      17'd49294: data = 8'hfd;
      17'd49295: data = 8'hfd;
      17'd49296: data = 8'hfe;
      17'd49297: data = 8'hfe;
      17'd49298: data = 8'h00;
      17'd49299: data = 8'h00;
      17'd49300: data = 8'h00;
      17'd49301: data = 8'h01;
      17'd49302: data = 8'h00;
      17'd49303: data = 8'h00;
      17'd49304: data = 8'hfe;
      17'd49305: data = 8'hfe;
      17'd49306: data = 8'hfd;
      17'd49307: data = 8'hfd;
      17'd49308: data = 8'hfd;
      17'd49309: data = 8'hfd;
      17'd49310: data = 8'hfe;
      17'd49311: data = 8'h00;
      17'd49312: data = 8'h00;
      17'd49313: data = 8'h00;
      17'd49314: data = 8'h00;
      17'd49315: data = 8'h00;
      17'd49316: data = 8'h00;
      17'd49317: data = 8'h00;
      17'd49318: data = 8'h00;
      17'd49319: data = 8'hfe;
      17'd49320: data = 8'h00;
      17'd49321: data = 8'hfe;
      17'd49322: data = 8'hfc;
      17'd49323: data = 8'hfd;
      17'd49324: data = 8'hfe;
      17'd49325: data = 8'hfd;
      17'd49326: data = 8'hfd;
      17'd49327: data = 8'h00;
      17'd49328: data = 8'h00;
      17'd49329: data = 8'h00;
      17'd49330: data = 8'h00;
      17'd49331: data = 8'h00;
      17'd49332: data = 8'h00;
      17'd49333: data = 8'h01;
      17'd49334: data = 8'h00;
      17'd49335: data = 8'hfe;
      17'd49336: data = 8'h00;
      17'd49337: data = 8'hfe;
      17'd49338: data = 8'hfd;
      17'd49339: data = 8'hfd;
      17'd49340: data = 8'hfe;
      17'd49341: data = 8'h00;
      17'd49342: data = 8'hfe;
      17'd49343: data = 8'hfd;
      17'd49344: data = 8'h00;
      17'd49345: data = 8'h01;
      17'd49346: data = 8'h01;
      17'd49347: data = 8'h00;
      17'd49348: data = 8'h00;
      17'd49349: data = 8'hfe;
      17'd49350: data = 8'hfe;
      17'd49351: data = 8'hfe;
      17'd49352: data = 8'hfd;
      17'd49353: data = 8'hfd;
      17'd49354: data = 8'hfd;
      17'd49355: data = 8'hfc;
      17'd49356: data = 8'hfd;
      17'd49357: data = 8'hfc;
      17'd49358: data = 8'hfe;
      17'd49359: data = 8'hfe;
      17'd49360: data = 8'h00;
      17'd49361: data = 8'h00;
      17'd49362: data = 8'h00;
      17'd49363: data = 8'h01;
      17'd49364: data = 8'h00;
      17'd49365: data = 8'hfe;
      17'd49366: data = 8'hfe;
      17'd49367: data = 8'hfe;
      17'd49368: data = 8'h00;
      17'd49369: data = 8'h01;
      17'd49370: data = 8'h00;
      17'd49371: data = 8'h00;
      17'd49372: data = 8'h00;
      17'd49373: data = 8'h00;
      17'd49374: data = 8'h00;
      17'd49375: data = 8'hfd;
      17'd49376: data = 8'hfd;
      17'd49377: data = 8'hfe;
      17'd49378: data = 8'hfe;
      17'd49379: data = 8'hfe;
      17'd49380: data = 8'h00;
      17'd49381: data = 8'hfe;
      17'd49382: data = 8'hfd;
      17'd49383: data = 8'hfe;
      17'd49384: data = 8'h00;
      17'd49385: data = 8'h00;
      17'd49386: data = 8'hfe;
      17'd49387: data = 8'h00;
      17'd49388: data = 8'hfe;
      17'd49389: data = 8'hfd;
      17'd49390: data = 8'hfe;
      17'd49391: data = 8'hfe;
      17'd49392: data = 8'hfe;
      17'd49393: data = 8'h00;
      17'd49394: data = 8'hfe;
      17'd49395: data = 8'hfe;
      17'd49396: data = 8'hfe;
      17'd49397: data = 8'hfe;
      17'd49398: data = 8'h00;
      17'd49399: data = 8'h00;
      17'd49400: data = 8'h00;
      17'd49401: data = 8'hfe;
      17'd49402: data = 8'h00;
      17'd49403: data = 8'h00;
      17'd49404: data = 8'h00;
      17'd49405: data = 8'h00;
      17'd49406: data = 8'h00;
      17'd49407: data = 8'hfe;
      17'd49408: data = 8'hfd;
      17'd49409: data = 8'hfe;
      17'd49410: data = 8'h00;
      17'd49411: data = 8'hfd;
      17'd49412: data = 8'hfe;
      17'd49413: data = 8'h00;
      17'd49414: data = 8'h00;
      17'd49415: data = 8'h00;
      17'd49416: data = 8'hfe;
      17'd49417: data = 8'h00;
      17'd49418: data = 8'hfe;
      17'd49419: data = 8'h01;
      17'd49420: data = 8'h00;
      17'd49421: data = 8'hfe;
      17'd49422: data = 8'h00;
      17'd49423: data = 8'hfe;
      17'd49424: data = 8'hfe;
      17'd49425: data = 8'h00;
      17'd49426: data = 8'hfe;
      17'd49427: data = 8'hfd;
      17'd49428: data = 8'hfe;
      17'd49429: data = 8'h00;
      17'd49430: data = 8'h00;
      17'd49431: data = 8'h01;
      17'd49432: data = 8'h01;
      17'd49433: data = 8'h00;
      17'd49434: data = 8'h01;
      17'd49435: data = 8'h01;
      17'd49436: data = 8'h01;
      17'd49437: data = 8'h01;
      17'd49438: data = 8'h00;
      17'd49439: data = 8'hfe;
      17'd49440: data = 8'h00;
      17'd49441: data = 8'hfe;
      17'd49442: data = 8'hfe;
      17'd49443: data = 8'h00;
      17'd49444: data = 8'h00;
      17'd49445: data = 8'h00;
      17'd49446: data = 8'h00;
      17'd49447: data = 8'h00;
      17'd49448: data = 8'h01;
      17'd49449: data = 8'h00;
      17'd49450: data = 8'h00;
      17'd49451: data = 8'h00;
      17'd49452: data = 8'hfe;
      17'd49453: data = 8'h00;
      17'd49454: data = 8'hfe;
      17'd49455: data = 8'hfe;
      17'd49456: data = 8'h00;
      17'd49457: data = 8'h00;
      17'd49458: data = 8'h01;
      17'd49459: data = 8'h01;
      17'd49460: data = 8'h01;
      17'd49461: data = 8'h01;
      17'd49462: data = 8'h00;
      17'd49463: data = 8'h01;
      17'd49464: data = 8'h00;
      17'd49465: data = 8'h00;
      17'd49466: data = 8'h00;
      17'd49467: data = 8'h00;
      17'd49468: data = 8'h00;
      17'd49469: data = 8'h00;
      17'd49470: data = 8'hfe;
      17'd49471: data = 8'hfd;
      17'd49472: data = 8'hfe;
      17'd49473: data = 8'h00;
      17'd49474: data = 8'h01;
      17'd49475: data = 8'h00;
      17'd49476: data = 8'h00;
      17'd49477: data = 8'h00;
      17'd49478: data = 8'h00;
      17'd49479: data = 8'h01;
      17'd49480: data = 8'hfe;
      17'd49481: data = 8'h00;
      17'd49482: data = 8'hfd;
      17'd49483: data = 8'hfe;
      17'd49484: data = 8'hfe;
      17'd49485: data = 8'h00;
      17'd49486: data = 8'hfe;
      17'd49487: data = 8'h00;
      17'd49488: data = 8'h00;
      17'd49489: data = 8'h01;
      17'd49490: data = 8'h01;
      17'd49491: data = 8'h01;
      17'd49492: data = 8'h01;
      17'd49493: data = 8'h00;
      17'd49494: data = 8'h01;
      17'd49495: data = 8'h00;
      17'd49496: data = 8'h00;
      17'd49497: data = 8'h00;
      17'd49498: data = 8'hfe;
      17'd49499: data = 8'h00;
      17'd49500: data = 8'hfe;
      17'd49501: data = 8'hfd;
      17'd49502: data = 8'hfe;
      17'd49503: data = 8'h00;
      17'd49504: data = 8'h00;
      17'd49505: data = 8'hfe;
      17'd49506: data = 8'hfe;
      17'd49507: data = 8'h00;
      17'd49508: data = 8'h01;
      17'd49509: data = 8'h02;
      17'd49510: data = 8'h02;
      17'd49511: data = 8'h00;
      17'd49512: data = 8'h00;
      17'd49513: data = 8'h01;
      17'd49514: data = 8'hfe;
      17'd49515: data = 8'hfe;
      17'd49516: data = 8'hfe;
      17'd49517: data = 8'hfd;
      17'd49518: data = 8'hfe;
      17'd49519: data = 8'h00;
      17'd49520: data = 8'h00;
      17'd49521: data = 8'h00;
      17'd49522: data = 8'h00;
      17'd49523: data = 8'h00;
      17'd49524: data = 8'h01;
      17'd49525: data = 8'h01;
      17'd49526: data = 8'h01;
      17'd49527: data = 8'h01;
      17'd49528: data = 8'hfe;
      17'd49529: data = 8'hfe;
      17'd49530: data = 8'hfe;
      17'd49531: data = 8'hfe;
      17'd49532: data = 8'hfd;
      17'd49533: data = 8'hfe;
      17'd49534: data = 8'h00;
      17'd49535: data = 8'hfd;
      17'd49536: data = 8'hfe;
      17'd49537: data = 8'h00;
      17'd49538: data = 8'h01;
      17'd49539: data = 8'h01;
      17'd49540: data = 8'h00;
      17'd49541: data = 8'h00;
      17'd49542: data = 8'h00;
      17'd49543: data = 8'h00;
      17'd49544: data = 8'hfe;
      17'd49545: data = 8'hfe;
      17'd49546: data = 8'h00;
      17'd49547: data = 8'h00;
      17'd49548: data = 8'hfd;
      17'd49549: data = 8'hfc;
      17'd49550: data = 8'hfe;
      17'd49551: data = 8'hfd;
      17'd49552: data = 8'hfe;
      17'd49553: data = 8'hfe;
      17'd49554: data = 8'hfe;
      17'd49555: data = 8'hfe;
      17'd49556: data = 8'hfe;
      17'd49557: data = 8'h00;
      17'd49558: data = 8'hfe;
      17'd49559: data = 8'hfe;
      17'd49560: data = 8'hfd;
      17'd49561: data = 8'hfc;
      17'd49562: data = 8'hfc;
      17'd49563: data = 8'hfd;
      17'd49564: data = 8'hfd;
      17'd49565: data = 8'hfc;
      17'd49566: data = 8'hfe;
      17'd49567: data = 8'hfe;
      17'd49568: data = 8'h00;
      17'd49569: data = 8'h01;
      17'd49570: data = 8'h00;
      17'd49571: data = 8'h00;
      17'd49572: data = 8'h00;
      17'd49573: data = 8'h00;
      17'd49574: data = 8'hfe;
      17'd49575: data = 8'hfe;
      17'd49576: data = 8'hfd;
      17'd49577: data = 8'hfd;
      17'd49578: data = 8'hfd;
      17'd49579: data = 8'hfc;
      17'd49580: data = 8'hfd;
      17'd49581: data = 8'hfe;
      17'd49582: data = 8'hfd;
      17'd49583: data = 8'hfd;
      17'd49584: data = 8'hfe;
      17'd49585: data = 8'hfe;
      17'd49586: data = 8'hfd;
      17'd49587: data = 8'hfe;
      17'd49588: data = 8'h00;
      17'd49589: data = 8'h00;
      17'd49590: data = 8'hfe;
      17'd49591: data = 8'hfe;
      17'd49592: data = 8'hfe;
      17'd49593: data = 8'hfd;
      17'd49594: data = 8'h00;
      17'd49595: data = 8'hfd;
      17'd49596: data = 8'hfe;
      17'd49597: data = 8'hfe;
      17'd49598: data = 8'hfe;
      17'd49599: data = 8'hfe;
      17'd49600: data = 8'hfd;
      17'd49601: data = 8'h00;
      17'd49602: data = 8'hfd;
      17'd49603: data = 8'h00;
      17'd49604: data = 8'h00;
      17'd49605: data = 8'h00;
      17'd49606: data = 8'hfe;
      17'd49607: data = 8'h00;
      17'd49608: data = 8'h00;
      17'd49609: data = 8'hfd;
      17'd49610: data = 8'hfe;
      17'd49611: data = 8'hfd;
      17'd49612: data = 8'hfd;
      17'd49613: data = 8'hfe;
      17'd49614: data = 8'hfe;
      17'd49615: data = 8'hfe;
      17'd49616: data = 8'hfe;
      17'd49617: data = 8'hfe;
      17'd49618: data = 8'h00;
      17'd49619: data = 8'h00;
      17'd49620: data = 8'h00;
      17'd49621: data = 8'h00;
      17'd49622: data = 8'h00;
      17'd49623: data = 8'hfe;
      17'd49624: data = 8'hfe;
      17'd49625: data = 8'hfe;
      17'd49626: data = 8'hfe;
      17'd49627: data = 8'hfd;
      17'd49628: data = 8'hfe;
      17'd49629: data = 8'hfe;
      17'd49630: data = 8'hfe;
      17'd49631: data = 8'hfe;
      17'd49632: data = 8'hfe;
      17'd49633: data = 8'h00;
      17'd49634: data = 8'h00;
      17'd49635: data = 8'h01;
      17'd49636: data = 8'h00;
      17'd49637: data = 8'hfe;
      17'd49638: data = 8'h00;
      17'd49639: data = 8'h01;
      17'd49640: data = 8'h00;
      17'd49641: data = 8'h00;
      17'd49642: data = 8'h00;
      17'd49643: data = 8'h00;
      17'd49644: data = 8'h00;
      17'd49645: data = 8'h00;
      17'd49646: data = 8'hfe;
      17'd49647: data = 8'hfe;
      17'd49648: data = 8'h01;
      17'd49649: data = 8'h00;
      17'd49650: data = 8'h01;
      17'd49651: data = 8'h01;
      17'd49652: data = 8'hfe;
      17'd49653: data = 8'h01;
      17'd49654: data = 8'h01;
      17'd49655: data = 8'h02;
      17'd49656: data = 8'h00;
      17'd49657: data = 8'h00;
      17'd49658: data = 8'h00;
      17'd49659: data = 8'h00;
      17'd49660: data = 8'h00;
      17'd49661: data = 8'hfd;
      17'd49662: data = 8'hfe;
      17'd49663: data = 8'hfe;
      17'd49664: data = 8'hfe;
      17'd49665: data = 8'hfe;
      17'd49666: data = 8'hfe;
      17'd49667: data = 8'h00;
      17'd49668: data = 8'h00;
      17'd49669: data = 8'h01;
      17'd49670: data = 8'h00;
      17'd49671: data = 8'h00;
      17'd49672: data = 8'h00;
      17'd49673: data = 8'h00;
      17'd49674: data = 8'h00;
      17'd49675: data = 8'h00;
      17'd49676: data = 8'hfe;
      17'd49677: data = 8'hfd;
      17'd49678: data = 8'hfe;
      17'd49679: data = 8'h00;
      17'd49680: data = 8'h01;
      17'd49681: data = 8'h00;
      17'd49682: data = 8'h00;
      17'd49683: data = 8'h00;
      17'd49684: data = 8'hfe;
      17'd49685: data = 8'h00;
      17'd49686: data = 8'h01;
      17'd49687: data = 8'h01;
      17'd49688: data = 8'h01;
      17'd49689: data = 8'h00;
      17'd49690: data = 8'h00;
      17'd49691: data = 8'h00;
      17'd49692: data = 8'h00;
      17'd49693: data = 8'h01;
      17'd49694: data = 8'h00;
      17'd49695: data = 8'h00;
      17'd49696: data = 8'h01;
      17'd49697: data = 8'h01;
      17'd49698: data = 8'h00;
      17'd49699: data = 8'h01;
      17'd49700: data = 8'h02;
      17'd49701: data = 8'h01;
      17'd49702: data = 8'h01;
      17'd49703: data = 8'h01;
      17'd49704: data = 8'h01;
      17'd49705: data = 8'h02;
      17'd49706: data = 8'h01;
      17'd49707: data = 8'h01;
      17'd49708: data = 8'h00;
      17'd49709: data = 8'h00;
      17'd49710: data = 8'hfe;
      17'd49711: data = 8'hfe;
      17'd49712: data = 8'hfe;
      17'd49713: data = 8'hfe;
      17'd49714: data = 8'h00;
      17'd49715: data = 8'hfe;
      17'd49716: data = 8'h00;
      17'd49717: data = 8'h00;
      17'd49718: data = 8'h01;
      17'd49719: data = 8'h01;
      17'd49720: data = 8'h00;
      17'd49721: data = 8'h00;
      17'd49722: data = 8'h00;
      17'd49723: data = 8'hfe;
      17'd49724: data = 8'hfd;
      17'd49725: data = 8'hfd;
      17'd49726: data = 8'hfe;
      17'd49727: data = 8'hfd;
      17'd49728: data = 8'hfd;
      17'd49729: data = 8'h00;
      17'd49730: data = 8'hfe;
      17'd49731: data = 8'h00;
      17'd49732: data = 8'h00;
      17'd49733: data = 8'h00;
      17'd49734: data = 8'h01;
      17'd49735: data = 8'h01;
      17'd49736: data = 8'h01;
      17'd49737: data = 8'h00;
      17'd49738: data = 8'h00;
      17'd49739: data = 8'h00;
      17'd49740: data = 8'hfe;
      17'd49741: data = 8'hfe;
      17'd49742: data = 8'hfe;
      17'd49743: data = 8'hfe;
      17'd49744: data = 8'h00;
      17'd49745: data = 8'h00;
      17'd49746: data = 8'h01;
      17'd49747: data = 8'h01;
      17'd49748: data = 8'h01;
      17'd49749: data = 8'h01;
      17'd49750: data = 8'h02;
      17'd49751: data = 8'h01;
      17'd49752: data = 8'h01;
      17'd49753: data = 8'h01;
      17'd49754: data = 8'hfe;
      17'd49755: data = 8'h00;
      17'd49756: data = 8'h00;
      17'd49757: data = 8'h00;
      17'd49758: data = 8'hfe;
      17'd49759: data = 8'hfe;
      17'd49760: data = 8'hfe;
      17'd49761: data = 8'hfe;
      17'd49762: data = 8'h00;
      17'd49763: data = 8'hfe;
      17'd49764: data = 8'h00;
      17'd49765: data = 8'h01;
      17'd49766: data = 8'h02;
      17'd49767: data = 8'h01;
      17'd49768: data = 8'h01;
      17'd49769: data = 8'h01;
      17'd49770: data = 8'h01;
      17'd49771: data = 8'h00;
      17'd49772: data = 8'h00;
      17'd49773: data = 8'h00;
      17'd49774: data = 8'hfe;
      17'd49775: data = 8'hfd;
      17'd49776: data = 8'hfe;
      17'd49777: data = 8'h00;
      17'd49778: data = 8'h00;
      17'd49779: data = 8'h02;
      17'd49780: data = 8'h02;
      17'd49781: data = 8'h01;
      17'd49782: data = 8'h00;
      17'd49783: data = 8'h00;
      17'd49784: data = 8'h00;
      17'd49785: data = 8'h00;
      17'd49786: data = 8'hfe;
      17'd49787: data = 8'hfe;
      17'd49788: data = 8'hfd;
      17'd49789: data = 8'hfd;
      17'd49790: data = 8'hfe;
      17'd49791: data = 8'hfd;
      17'd49792: data = 8'hfd;
      17'd49793: data = 8'hfe;
      17'd49794: data = 8'h00;
      17'd49795: data = 8'h00;
      17'd49796: data = 8'h00;
      17'd49797: data = 8'h00;
      17'd49798: data = 8'h00;
      17'd49799: data = 8'h00;
      17'd49800: data = 8'h00;
      17'd49801: data = 8'hfe;
      17'd49802: data = 8'hfe;
      17'd49803: data = 8'hfe;
      17'd49804: data = 8'hfe;
      17'd49805: data = 8'h00;
      17'd49806: data = 8'hfe;
      17'd49807: data = 8'hfe;
      17'd49808: data = 8'hfe;
      17'd49809: data = 8'hfe;
      17'd49810: data = 8'h00;
      17'd49811: data = 8'h00;
      17'd49812: data = 8'h00;
      17'd49813: data = 8'hfe;
      17'd49814: data = 8'hfe;
      17'd49815: data = 8'hfe;
      17'd49816: data = 8'hfe;
      17'd49817: data = 8'hfe;
      17'd49818: data = 8'hfd;
      17'd49819: data = 8'hfe;
      17'd49820: data = 8'hfe;
      17'd49821: data = 8'hfe;
      17'd49822: data = 8'hfe;
      17'd49823: data = 8'hfe;
      17'd49824: data = 8'hfe;
      17'd49825: data = 8'hfe;
      17'd49826: data = 8'hfe;
      17'd49827: data = 8'hfe;
      17'd49828: data = 8'hfe;
      17'd49829: data = 8'hfe;
      17'd49830: data = 8'hfe;
      17'd49831: data = 8'hfe;
      17'd49832: data = 8'hfe;
      17'd49833: data = 8'h00;
      17'd49834: data = 8'h00;
      17'd49835: data = 8'hfe;
      17'd49836: data = 8'hfe;
      17'd49837: data = 8'h00;
      17'd49838: data = 8'h00;
      17'd49839: data = 8'hfe;
      17'd49840: data = 8'hfe;
      17'd49841: data = 8'hfe;
      17'd49842: data = 8'hfe;
      17'd49843: data = 8'hfe;
      17'd49844: data = 8'hfe;
      17'd49845: data = 8'hfe;
      17'd49846: data = 8'hfd;
      17'd49847: data = 8'hfd;
      17'd49848: data = 8'hfd;
      17'd49849: data = 8'h00;
      17'd49850: data = 8'hfe;
      17'd49851: data = 8'hfe;
      17'd49852: data = 8'hfe;
      17'd49853: data = 8'hfe;
      17'd49854: data = 8'h00;
      17'd49855: data = 8'hfe;
      17'd49856: data = 8'hfe;
      17'd49857: data = 8'h00;
      17'd49858: data = 8'hfe;
      17'd49859: data = 8'hfe;
      17'd49860: data = 8'hfe;
      17'd49861: data = 8'hfd;
      17'd49862: data = 8'hfd;
      17'd49863: data = 8'hfd;
      17'd49864: data = 8'hfe;
      17'd49865: data = 8'hfe;
      17'd49866: data = 8'hfe;
      17'd49867: data = 8'h00;
      17'd49868: data = 8'h00;
      17'd49869: data = 8'h00;
      17'd49870: data = 8'h00;
      17'd49871: data = 8'h00;
      17'd49872: data = 8'hfe;
      17'd49873: data = 8'hfe;
      17'd49874: data = 8'hfe;
      17'd49875: data = 8'hfe;
      17'd49876: data = 8'hfd;
      17'd49877: data = 8'hfd;
      17'd49878: data = 8'hfe;
      17'd49879: data = 8'h00;
      17'd49880: data = 8'h00;
      17'd49881: data = 8'h00;
      17'd49882: data = 8'h02;
      17'd49883: data = 8'h01;
      17'd49884: data = 8'h01;
      17'd49885: data = 8'h01;
      17'd49886: data = 8'hfe;
      17'd49887: data = 8'hfe;
      17'd49888: data = 8'hfd;
      17'd49889: data = 8'hfd;
      17'd49890: data = 8'hfd;
      17'd49891: data = 8'hfd;
      17'd49892: data = 8'hfd;
      17'd49893: data = 8'h00;
      17'd49894: data = 8'h01;
      17'd49895: data = 8'h00;
      17'd49896: data = 8'h01;
      17'd49897: data = 8'h02;
      17'd49898: data = 8'h02;
      17'd49899: data = 8'h01;
      17'd49900: data = 8'h01;
      17'd49901: data = 8'h00;
      17'd49902: data = 8'hfe;
      17'd49903: data = 8'hfd;
      17'd49904: data = 8'hfd;
      17'd49905: data = 8'hfe;
      17'd49906: data = 8'hfd;
      17'd49907: data = 8'hfe;
      17'd49908: data = 8'h00;
      17'd49909: data = 8'h00;
      17'd49910: data = 8'h01;
      17'd49911: data = 8'h02;
      17'd49912: data = 8'h01;
      17'd49913: data = 8'h02;
      17'd49914: data = 8'h02;
      17'd49915: data = 8'h01;
      17'd49916: data = 8'hfe;
      17'd49917: data = 8'hfe;
      17'd49918: data = 8'hfd;
      17'd49919: data = 8'hfd;
      17'd49920: data = 8'hfd;
      17'd49921: data = 8'hfd;
      17'd49922: data = 8'hfd;
      17'd49923: data = 8'hfe;
      17'd49924: data = 8'h00;
      17'd49925: data = 8'h02;
      17'd49926: data = 8'h01;
      17'd49927: data = 8'h00;
      17'd49928: data = 8'h01;
      17'd49929: data = 8'h01;
      17'd49930: data = 8'hfe;
      17'd49931: data = 8'hfe;
      17'd49932: data = 8'hfe;
      17'd49933: data = 8'hfd;
      17'd49934: data = 8'hfe;
      17'd49935: data = 8'hfe;
      17'd49936: data = 8'h00;
      17'd49937: data = 8'h01;
      17'd49938: data = 8'h02;
      17'd49939: data = 8'h04;
      17'd49940: data = 8'h04;
      17'd49941: data = 8'h02;
      17'd49942: data = 8'h01;
      17'd49943: data = 8'h02;
      17'd49944: data = 8'h01;
      17'd49945: data = 8'h00;
      17'd49946: data = 8'h00;
      17'd49947: data = 8'hfe;
      17'd49948: data = 8'h00;
      17'd49949: data = 8'h00;
      17'd49950: data = 8'h00;
      17'd49951: data = 8'hfe;
      17'd49952: data = 8'h01;
      17'd49953: data = 8'h02;
      17'd49954: data = 8'h02;
      17'd49955: data = 8'h02;
      17'd49956: data = 8'h01;
      17'd49957: data = 8'h01;
      17'd49958: data = 8'h01;
      17'd49959: data = 8'h01;
      17'd49960: data = 8'h00;
      17'd49961: data = 8'hfe;
      17'd49962: data = 8'hfe;
      17'd49963: data = 8'h00;
      17'd49964: data = 8'h01;
      17'd49965: data = 8'h01;
      17'd49966: data = 8'h00;
      17'd49967: data = 8'h02;
      17'd49968: data = 8'h01;
      17'd49969: data = 8'h00;
      17'd49970: data = 8'h01;
      17'd49971: data = 8'h00;
      17'd49972: data = 8'h00;
      17'd49973: data = 8'hfe;
      17'd49974: data = 8'hfe;
      17'd49975: data = 8'hfe;
      17'd49976: data = 8'hfe;
      17'd49977: data = 8'hfd;
      17'd49978: data = 8'hfd;
      17'd49979: data = 8'h00;
      17'd49980: data = 8'h00;
      17'd49981: data = 8'h00;
      17'd49982: data = 8'h01;
      17'd49983: data = 8'h01;
      17'd49984: data = 8'h01;
      17'd49985: data = 8'h01;
      17'd49986: data = 8'h00;
      17'd49987: data = 8'hfe;
      17'd49988: data = 8'hfe;
      17'd49989: data = 8'hfd;
      17'd49990: data = 8'hfc;
      17'd49991: data = 8'hfd;
      17'd49992: data = 8'hfd;
      17'd49993: data = 8'hfe;
      17'd49994: data = 8'hfe;
      17'd49995: data = 8'hfe;
      17'd49996: data = 8'h01;
      17'd49997: data = 8'h01;
      17'd49998: data = 8'h00;
      17'd49999: data = 8'h02;
      17'd50000: data = 8'h01;
      17'd50001: data = 8'hfe;
      17'd50002: data = 8'h00;
      17'd50003: data = 8'hfe;
      17'd50004: data = 8'hfd;
      17'd50005: data = 8'hfe;
      17'd50006: data = 8'hfd;
      17'd50007: data = 8'hfd;
      17'd50008: data = 8'hfe;
      17'd50009: data = 8'h00;
      17'd50010: data = 8'hfe;
      17'd50011: data = 8'h01;
      17'd50012: data = 8'h01;
      17'd50013: data = 8'h00;
      17'd50014: data = 8'h00;
      17'd50015: data = 8'hfe;
      17'd50016: data = 8'hfd;
      17'd50017: data = 8'hfd;
      17'd50018: data = 8'hfd;
      17'd50019: data = 8'hfc;
      17'd50020: data = 8'hfd;
      17'd50021: data = 8'hfe;
      17'd50022: data = 8'hfd;
      17'd50023: data = 8'h00;
      17'd50024: data = 8'h01;
      17'd50025: data = 8'h01;
      17'd50026: data = 8'h01;
      17'd50027: data = 8'h00;
      17'd50028: data = 8'hfe;
      17'd50029: data = 8'hfd;
      17'd50030: data = 8'hfd;
      17'd50031: data = 8'hfe;
      17'd50032: data = 8'hfc;
      17'd50033: data = 8'hfc;
      17'd50034: data = 8'hfc;
      17'd50035: data = 8'hfd;
      17'd50036: data = 8'hfe;
      17'd50037: data = 8'hfe;
      17'd50038: data = 8'hfe;
      17'd50039: data = 8'h00;
      17'd50040: data = 8'h00;
      17'd50041: data = 8'h00;
      17'd50042: data = 8'hfe;
      17'd50043: data = 8'hfe;
      17'd50044: data = 8'hfe;
      17'd50045: data = 8'hfe;
      17'd50046: data = 8'hfe;
      17'd50047: data = 8'hfc;
      17'd50048: data = 8'hfc;
      17'd50049: data = 8'hfe;
      17'd50050: data = 8'hfe;
      17'd50051: data = 8'hfe;
      17'd50052: data = 8'h00;
      17'd50053: data = 8'h01;
      17'd50054: data = 8'h01;
      17'd50055: data = 8'h01;
      17'd50056: data = 8'h01;
      17'd50057: data = 8'h00;
      17'd50058: data = 8'hfe;
      17'd50059: data = 8'hfd;
      17'd50060: data = 8'hfd;
      17'd50061: data = 8'hfd;
      17'd50062: data = 8'hfd;
      17'd50063: data = 8'hfd;
      17'd50064: data = 8'hfe;
      17'd50065: data = 8'h00;
      17'd50066: data = 8'h00;
      17'd50067: data = 8'h01;
      17'd50068: data = 8'h01;
      17'd50069: data = 8'h01;
      17'd50070: data = 8'h02;
      17'd50071: data = 8'h01;
      17'd50072: data = 8'h00;
      17'd50073: data = 8'h00;
      17'd50074: data = 8'hfe;
      17'd50075: data = 8'hfc;
      17'd50076: data = 8'hfd;
      17'd50077: data = 8'hfd;
      17'd50078: data = 8'hfd;
      17'd50079: data = 8'hfe;
      17'd50080: data = 8'hfe;
      17'd50081: data = 8'h00;
      17'd50082: data = 8'hfe;
      17'd50083: data = 8'h00;
      17'd50084: data = 8'h01;
      17'd50085: data = 8'hfe;
      17'd50086: data = 8'hfe;
      17'd50087: data = 8'hfe;
      17'd50088: data = 8'hfe;
      17'd50089: data = 8'hfd;
      17'd50090: data = 8'hfd;
      17'd50091: data = 8'hfd;
      17'd50092: data = 8'hfd;
      17'd50093: data = 8'hfe;
      17'd50094: data = 8'hfe;
      17'd50095: data = 8'hfe;
      17'd50096: data = 8'h00;
      17'd50097: data = 8'h00;
      17'd50098: data = 8'h00;
      17'd50099: data = 8'h00;
      17'd50100: data = 8'h00;
      17'd50101: data = 8'hfe;
      17'd50102: data = 8'h00;
      17'd50103: data = 8'h00;
      17'd50104: data = 8'h00;
      17'd50105: data = 8'hfe;
      17'd50106: data = 8'hfd;
      17'd50107: data = 8'hfd;
      17'd50108: data = 8'hfd;
      17'd50109: data = 8'h00;
      17'd50110: data = 8'h01;
      17'd50111: data = 8'h01;
      17'd50112: data = 8'h01;
      17'd50113: data = 8'h01;
      17'd50114: data = 8'h01;
      17'd50115: data = 8'h00;
      17'd50116: data = 8'h00;
      17'd50117: data = 8'hfe;
      17'd50118: data = 8'hfe;
      17'd50119: data = 8'hfe;
      17'd50120: data = 8'h00;
      17'd50121: data = 8'h00;
      17'd50122: data = 8'h00;
      17'd50123: data = 8'hfe;
      17'd50124: data = 8'hfe;
      17'd50125: data = 8'h00;
      17'd50126: data = 8'h01;
      17'd50127: data = 8'h00;
      17'd50128: data = 8'h00;
      17'd50129: data = 8'h00;
      17'd50130: data = 8'hfe;
      17'd50131: data = 8'h00;
      17'd50132: data = 8'h00;
      17'd50133: data = 8'hfe;
      17'd50134: data = 8'h00;
      17'd50135: data = 8'h00;
      17'd50136: data = 8'h01;
      17'd50137: data = 8'h01;
      17'd50138: data = 8'hfe;
      17'd50139: data = 8'hfe;
      17'd50140: data = 8'h00;
      17'd50141: data = 8'h00;
      17'd50142: data = 8'hfe;
      17'd50143: data = 8'hfe;
      17'd50144: data = 8'hfe;
      17'd50145: data = 8'hfd;
      17'd50146: data = 8'hfd;
      17'd50147: data = 8'hfe;
      17'd50148: data = 8'hfe;
      17'd50149: data = 8'h00;
      17'd50150: data = 8'h01;
      17'd50151: data = 8'h01;
      17'd50152: data = 8'h00;
      17'd50153: data = 8'h01;
      17'd50154: data = 8'h00;
      17'd50155: data = 8'h00;
      17'd50156: data = 8'h00;
      17'd50157: data = 8'hfe;
      17'd50158: data = 8'hfe;
      17'd50159: data = 8'hfe;
      17'd50160: data = 8'h00;
      17'd50161: data = 8'hfe;
      17'd50162: data = 8'hfe;
      17'd50163: data = 8'hfe;
      17'd50164: data = 8'h00;
      17'd50165: data = 8'h02;
      17'd50166: data = 8'h02;
      17'd50167: data = 8'h01;
      17'd50168: data = 8'h01;
      17'd50169: data = 8'h01;
      17'd50170: data = 8'h01;
      17'd50171: data = 8'h00;
      17'd50172: data = 8'hfe;
      17'd50173: data = 8'hfe;
      17'd50174: data = 8'hfe;
      17'd50175: data = 8'hfe;
      17'd50176: data = 8'hfd;
      17'd50177: data = 8'hfd;
      17'd50178: data = 8'h00;
      17'd50179: data = 8'h01;
      17'd50180: data = 8'h00;
      17'd50181: data = 8'h00;
      17'd50182: data = 8'h01;
      17'd50183: data = 8'h01;
      17'd50184: data = 8'h01;
      17'd50185: data = 8'h00;
      17'd50186: data = 8'h00;
      17'd50187: data = 8'hfe;
      17'd50188: data = 8'hfe;
      17'd50189: data = 8'hfd;
      17'd50190: data = 8'hfe;
      17'd50191: data = 8'hfe;
      17'd50192: data = 8'hfe;
      17'd50193: data = 8'h00;
      17'd50194: data = 8'h01;
      17'd50195: data = 8'h01;
      17'd50196: data = 8'h01;
      17'd50197: data = 8'h02;
      17'd50198: data = 8'h02;
      17'd50199: data = 8'h01;
      17'd50200: data = 8'h00;
      17'd50201: data = 8'h00;
      17'd50202: data = 8'hfe;
      17'd50203: data = 8'hfe;
      17'd50204: data = 8'hfe;
      17'd50205: data = 8'hfe;
      17'd50206: data = 8'hfe;
      17'd50207: data = 8'hfe;
      17'd50208: data = 8'h00;
      17'd50209: data = 8'h00;
      17'd50210: data = 8'h00;
      17'd50211: data = 8'h00;
      17'd50212: data = 8'h00;
      17'd50213: data = 8'h00;
      17'd50214: data = 8'h00;
      17'd50215: data = 8'h00;
      17'd50216: data = 8'hfe;
      17'd50217: data = 8'hfe;
      17'd50218: data = 8'hfd;
      17'd50219: data = 8'hfd;
      17'd50220: data = 8'hfe;
      17'd50221: data = 8'hfe;
      17'd50222: data = 8'hfe;
      17'd50223: data = 8'hfe;
      17'd50224: data = 8'h01;
      17'd50225: data = 8'h01;
      17'd50226: data = 8'h01;
      17'd50227: data = 8'h00;
      17'd50228: data = 8'h00;
      17'd50229: data = 8'h01;
      17'd50230: data = 8'h00;
      17'd50231: data = 8'hfd;
      17'd50232: data = 8'hfd;
      17'd50233: data = 8'hfd;
      17'd50234: data = 8'hfd;
      17'd50235: data = 8'hfd;
      17'd50236: data = 8'hfc;
      17'd50237: data = 8'hfe;
      17'd50238: data = 8'hfe;
      17'd50239: data = 8'hfe;
      17'd50240: data = 8'h00;
      17'd50241: data = 8'h00;
      17'd50242: data = 8'h00;
      17'd50243: data = 8'h00;
      17'd50244: data = 8'hfd;
      17'd50245: data = 8'hfd;
      17'd50246: data = 8'hfd;
      17'd50247: data = 8'hfd;
      17'd50248: data = 8'hfd;
      17'd50249: data = 8'hfd;
      17'd50250: data = 8'hfc;
      17'd50251: data = 8'hfd;
      17'd50252: data = 8'hfe;
      17'd50253: data = 8'h00;
      17'd50254: data = 8'h00;
      17'd50255: data = 8'h00;
      17'd50256: data = 8'h00;
      17'd50257: data = 8'h00;
      17'd50258: data = 8'hfe;
      17'd50259: data = 8'hfe;
      17'd50260: data = 8'hfe;
      17'd50261: data = 8'hfd;
      17'd50262: data = 8'hfe;
      17'd50263: data = 8'hfe;
      17'd50264: data = 8'hfe;
      17'd50265: data = 8'hfd;
      17'd50266: data = 8'h00;
      17'd50267: data = 8'h00;
      17'd50268: data = 8'h00;
      17'd50269: data = 8'h01;
      17'd50270: data = 8'h00;
      17'd50271: data = 8'h00;
      17'd50272: data = 8'hfe;
      17'd50273: data = 8'hfe;
      17'd50274: data = 8'hfd;
      17'd50275: data = 8'hfd;
      17'd50276: data = 8'hfe;
      17'd50277: data = 8'hfe;
      17'd50278: data = 8'hfe;
      17'd50279: data = 8'hfe;
      17'd50280: data = 8'h00;
      17'd50281: data = 8'hfe;
      17'd50282: data = 8'h00;
      17'd50283: data = 8'h01;
      17'd50284: data = 8'h01;
      17'd50285: data = 8'h01;
      17'd50286: data = 8'h01;
      17'd50287: data = 8'h01;
      17'd50288: data = 8'hfe;
      17'd50289: data = 8'hfe;
      17'd50290: data = 8'h00;
      17'd50291: data = 8'hfe;
      17'd50292: data = 8'h00;
      17'd50293: data = 8'hfe;
      17'd50294: data = 8'hfe;
      17'd50295: data = 8'h00;
      17'd50296: data = 8'h01;
      17'd50297: data = 8'h04;
      17'd50298: data = 8'h01;
      17'd50299: data = 8'h00;
      17'd50300: data = 8'h00;
      17'd50301: data = 8'h00;
      17'd50302: data = 8'hfe;
      17'd50303: data = 8'hfe;
      17'd50304: data = 8'hfe;
      17'd50305: data = 8'hfd;
      17'd50306: data = 8'hfe;
      17'd50307: data = 8'hfe;
      17'd50308: data = 8'hfd;
      17'd50309: data = 8'hfe;
      17'd50310: data = 8'hfe;
      17'd50311: data = 8'hfe;
      17'd50312: data = 8'h00;
      17'd50313: data = 8'h01;
      17'd50314: data = 8'h00;
      17'd50315: data = 8'h00;
      17'd50316: data = 8'h01;
      17'd50317: data = 8'h00;
      17'd50318: data = 8'h00;
      17'd50319: data = 8'h00;
      17'd50320: data = 8'hfe;
      17'd50321: data = 8'hfe;
      17'd50322: data = 8'h00;
      17'd50323: data = 8'hfe;
      17'd50324: data = 8'hfd;
      17'd50325: data = 8'h00;
      17'd50326: data = 8'h00;
      17'd50327: data = 8'h01;
      17'd50328: data = 8'h01;
      17'd50329: data = 8'h01;
      17'd50330: data = 8'h01;
      17'd50331: data = 8'h01;
      17'd50332: data = 8'h01;
      17'd50333: data = 8'hfe;
      17'd50334: data = 8'hfe;
      17'd50335: data = 8'hfe;
      17'd50336: data = 8'hfe;
      17'd50337: data = 8'hfd;
      17'd50338: data = 8'hfd;
      17'd50339: data = 8'hfd;
      17'd50340: data = 8'hfe;
      17'd50341: data = 8'hfe;
      17'd50342: data = 8'h00;
      17'd50343: data = 8'h00;
      17'd50344: data = 8'h00;
      17'd50345: data = 8'h00;
      17'd50346: data = 8'hfe;
      17'd50347: data = 8'h00;
      17'd50348: data = 8'hfe;
      17'd50349: data = 8'hfe;
      17'd50350: data = 8'hfe;
      17'd50351: data = 8'hfe;
      17'd50352: data = 8'hfe;
      17'd50353: data = 8'hfe;
      17'd50354: data = 8'hfe;
      17'd50355: data = 8'hfe;
      17'd50356: data = 8'h00;
      17'd50357: data = 8'h00;
      17'd50358: data = 8'h01;
      17'd50359: data = 8'h01;
      17'd50360: data = 8'h00;
      17'd50361: data = 8'h00;
      17'd50362: data = 8'h00;
      17'd50363: data = 8'h00;
      17'd50364: data = 8'hfe;
      17'd50365: data = 8'h00;
      17'd50366: data = 8'hfe;
      17'd50367: data = 8'hfe;
      17'd50368: data = 8'hfe;
      17'd50369: data = 8'hfe;
      17'd50370: data = 8'hfe;
      17'd50371: data = 8'h00;
      17'd50372: data = 8'h00;
      17'd50373: data = 8'h01;
      17'd50374: data = 8'h00;
      17'd50375: data = 8'h00;
      17'd50376: data = 8'h00;
      17'd50377: data = 8'h00;
      17'd50378: data = 8'h00;
      17'd50379: data = 8'h00;
      17'd50380: data = 8'h01;
      17'd50381: data = 8'hfe;
      17'd50382: data = 8'hfe;
      17'd50383: data = 8'h00;
      17'd50384: data = 8'h00;
      17'd50385: data = 8'h00;
      17'd50386: data = 8'h01;
      17'd50387: data = 8'h01;
      17'd50388: data = 8'h00;
      17'd50389: data = 8'h00;
      17'd50390: data = 8'h00;
      17'd50391: data = 8'h01;
      17'd50392: data = 8'hfe;
      17'd50393: data = 8'h00;
      17'd50394: data = 8'h00;
      17'd50395: data = 8'hfe;
      17'd50396: data = 8'hfe;
      17'd50397: data = 8'hfe;
      17'd50398: data = 8'hfe;
      17'd50399: data = 8'hfe;
      17'd50400: data = 8'h00;
      17'd50401: data = 8'h00;
      17'd50402: data = 8'h00;
      17'd50403: data = 8'h00;
      17'd50404: data = 8'h00;
      17'd50405: data = 8'h01;
      17'd50406: data = 8'hfe;
      17'd50407: data = 8'hfe;
      17'd50408: data = 8'hfe;
      17'd50409: data = 8'hfe;
      17'd50410: data = 8'hfe;
      17'd50411: data = 8'hfd;
      17'd50412: data = 8'hfe;
      17'd50413: data = 8'hfe;
      17'd50414: data = 8'h00;
      17'd50415: data = 8'h01;
      17'd50416: data = 8'h00;
      17'd50417: data = 8'h00;
      17'd50418: data = 8'h01;
      17'd50419: data = 8'h00;
      17'd50420: data = 8'h00;
      17'd50421: data = 8'hfe;
      17'd50422: data = 8'hfe;
      17'd50423: data = 8'h00;
      17'd50424: data = 8'h00;
      17'd50425: data = 8'h00;
      17'd50426: data = 8'h00;
      17'd50427: data = 8'h00;
      17'd50428: data = 8'h02;
      17'd50429: data = 8'h02;
      17'd50430: data = 8'h01;
      17'd50431: data = 8'h02;
      17'd50432: data = 8'h01;
      17'd50433: data = 8'h01;
      17'd50434: data = 8'h01;
      17'd50435: data = 8'h01;
      17'd50436: data = 8'h00;
      17'd50437: data = 8'h00;
      17'd50438: data = 8'h00;
      17'd50439: data = 8'h00;
      17'd50440: data = 8'hfe;
      17'd50441: data = 8'h00;
      17'd50442: data = 8'h01;
      17'd50443: data = 8'h01;
      17'd50444: data = 8'h00;
      17'd50445: data = 8'h01;
      17'd50446: data = 8'h02;
      17'd50447: data = 8'h02;
      17'd50448: data = 8'h01;
      17'd50449: data = 8'h00;
      17'd50450: data = 8'h01;
      17'd50451: data = 8'h00;
      17'd50452: data = 8'h00;
      17'd50453: data = 8'h00;
      17'd50454: data = 8'h00;
      17'd50455: data = 8'h00;
      17'd50456: data = 8'h00;
      17'd50457: data = 8'hfe;
      17'd50458: data = 8'h01;
      17'd50459: data = 8'h02;
      17'd50460: data = 8'h01;
      17'd50461: data = 8'h00;
      17'd50462: data = 8'h00;
      17'd50463: data = 8'h01;
      17'd50464: data = 8'h00;
      17'd50465: data = 8'hfe;
      17'd50466: data = 8'hfe;
      17'd50467: data = 8'hfe;
      17'd50468: data = 8'hfe;
      17'd50469: data = 8'hfd;
      17'd50470: data = 8'hfe;
      17'd50471: data = 8'hfe;
      17'd50472: data = 8'hfe;
      17'd50473: data = 8'h00;
      17'd50474: data = 8'h00;
      17'd50475: data = 8'h00;
      17'd50476: data = 8'h01;
      17'd50477: data = 8'h01;
      17'd50478: data = 8'h00;
      17'd50479: data = 8'h00;
      17'd50480: data = 8'h00;
      17'd50481: data = 8'hfe;
      17'd50482: data = 8'hfd;
      17'd50483: data = 8'hfd;
      17'd50484: data = 8'hfd;
      17'd50485: data = 8'hfd;
      17'd50486: data = 8'h00;
      17'd50487: data = 8'hfe;
      17'd50488: data = 8'h00;
      17'd50489: data = 8'hfe;
      17'd50490: data = 8'h00;
      17'd50491: data = 8'h02;
      17'd50492: data = 8'h00;
      17'd50493: data = 8'h00;
      17'd50494: data = 8'hfe;
      17'd50495: data = 8'hfe;
      17'd50496: data = 8'h00;
      17'd50497: data = 8'h00;
      17'd50498: data = 8'hfe;
      17'd50499: data = 8'h00;
      17'd50500: data = 8'h00;
      17'd50501: data = 8'hfe;
      17'd50502: data = 8'h00;
      17'd50503: data = 8'h00;
      17'd50504: data = 8'hfe;
      17'd50505: data = 8'h00;
      17'd50506: data = 8'hfe;
      17'd50507: data = 8'h00;
      17'd50508: data = 8'h01;
      17'd50509: data = 8'h00;
      17'd50510: data = 8'h00;
      17'd50511: data = 8'hfe;
      17'd50512: data = 8'hfe;
      17'd50513: data = 8'h00;
      17'd50514: data = 8'h00;
      17'd50515: data = 8'h00;
      17'd50516: data = 8'h00;
      17'd50517: data = 8'hfe;
      17'd50518: data = 8'hfe;
      17'd50519: data = 8'hfd;
      17'd50520: data = 8'h00;
      17'd50521: data = 8'h00;
      17'd50522: data = 8'hfe;
      17'd50523: data = 8'h01;
      17'd50524: data = 8'h00;
      17'd50525: data = 8'h00;
      17'd50526: data = 8'hfe;
      17'd50527: data = 8'hfe;
      17'd50528: data = 8'hfe;
      17'd50529: data = 8'hfe;
      17'd50530: data = 8'hfe;
      17'd50531: data = 8'hfd;
      17'd50532: data = 8'h00;
      17'd50533: data = 8'hfd;
      17'd50534: data = 8'h00;
      17'd50535: data = 8'h00;
      17'd50536: data = 8'hfe;
      17'd50537: data = 8'h00;
      17'd50538: data = 8'h00;
      17'd50539: data = 8'h00;
      17'd50540: data = 8'h00;
      17'd50541: data = 8'h00;
      17'd50542: data = 8'hfe;
      17'd50543: data = 8'h00;
      17'd50544: data = 8'h00;
      17'd50545: data = 8'hfe;
      17'd50546: data = 8'h00;
      17'd50547: data = 8'hfd;
      17'd50548: data = 8'hfe;
      17'd50549: data = 8'h00;
      17'd50550: data = 8'h00;
      17'd50551: data = 8'h00;
      17'd50552: data = 8'h00;
      17'd50553: data = 8'h02;
      17'd50554: data = 8'h01;
      17'd50555: data = 8'h00;
      17'd50556: data = 8'h00;
      17'd50557: data = 8'hfe;
      17'd50558: data = 8'h00;
      17'd50559: data = 8'hfe;
      17'd50560: data = 8'hfd;
      17'd50561: data = 8'hfe;
      17'd50562: data = 8'hfd;
      17'd50563: data = 8'hfe;
      17'd50564: data = 8'hfe;
      17'd50565: data = 8'hfe;
      17'd50566: data = 8'hfe;
      17'd50567: data = 8'hfe;
      17'd50568: data = 8'h00;
      17'd50569: data = 8'h01;
      17'd50570: data = 8'h01;
      17'd50571: data = 8'h01;
      17'd50572: data = 8'h01;
      17'd50573: data = 8'h00;
      17'd50574: data = 8'h00;
      17'd50575: data = 8'h01;
      17'd50576: data = 8'h00;
      17'd50577: data = 8'h00;
      17'd50578: data = 8'hfe;
      17'd50579: data = 8'h00;
      17'd50580: data = 8'h00;
      17'd50581: data = 8'h00;
      17'd50582: data = 8'hfe;
      17'd50583: data = 8'h00;
      17'd50584: data = 8'h01;
      17'd50585: data = 8'h00;
      17'd50586: data = 8'h00;
      17'd50587: data = 8'h01;
      17'd50588: data = 8'h00;
      17'd50589: data = 8'hfe;
      17'd50590: data = 8'hfe;
      17'd50591: data = 8'hfe;
      17'd50592: data = 8'hfe;
      17'd50593: data = 8'h00;
      17'd50594: data = 8'h00;
      17'd50595: data = 8'hfe;
      17'd50596: data = 8'hfe;
      17'd50597: data = 8'hfe;
      17'd50598: data = 8'h00;
      17'd50599: data = 8'hfe;
      17'd50600: data = 8'h00;
      17'd50601: data = 8'h01;
      17'd50602: data = 8'h01;
      17'd50603: data = 8'h00;
      17'd50604: data = 8'h00;
      17'd50605: data = 8'h00;
      17'd50606: data = 8'h00;
      17'd50607: data = 8'hfe;
      17'd50608: data = 8'hfe;
      17'd50609: data = 8'hfe;
      17'd50610: data = 8'hfe;
      17'd50611: data = 8'hfe;
      17'd50612: data = 8'h00;
      17'd50613: data = 8'h00;
      17'd50614: data = 8'h00;
      17'd50615: data = 8'h01;
      17'd50616: data = 8'h01;
      17'd50617: data = 8'h02;
      17'd50618: data = 8'h02;
      17'd50619: data = 8'h01;
      17'd50620: data = 8'h01;
      17'd50621: data = 8'h00;
      17'd50622: data = 8'h01;
      17'd50623: data = 8'h00;
      17'd50624: data = 8'hfd;
      17'd50625: data = 8'hfe;
      17'd50626: data = 8'hfe;
      17'd50627: data = 8'hfe;
      17'd50628: data = 8'hfe;
      17'd50629: data = 8'h00;
      17'd50630: data = 8'h00;
      17'd50631: data = 8'h00;
      17'd50632: data = 8'h01;
      17'd50633: data = 8'h00;
      17'd50634: data = 8'h00;
      17'd50635: data = 8'h00;
      17'd50636: data = 8'hfe;
      17'd50637: data = 8'h00;
      17'd50638: data = 8'h00;
      17'd50639: data = 8'h00;
      17'd50640: data = 8'hfe;
      17'd50641: data = 8'hfe;
      17'd50642: data = 8'hfe;
      17'd50643: data = 8'hfe;
      17'd50644: data = 8'h00;
      17'd50645: data = 8'hfe;
      17'd50646: data = 8'h00;
      17'd50647: data = 8'h00;
      17'd50648: data = 8'h00;
      17'd50649: data = 8'h01;
      17'd50650: data = 8'h01;
      17'd50651: data = 8'h01;
      17'd50652: data = 8'h01;
      17'd50653: data = 8'h02;
      17'd50654: data = 8'h00;
      17'd50655: data = 8'h00;
      17'd50656: data = 8'hfe;
      17'd50657: data = 8'hfe;
      17'd50658: data = 8'hfe;
      17'd50659: data = 8'hfd;
      17'd50660: data = 8'hfe;
      17'd50661: data = 8'hfe;
      17'd50662: data = 8'h00;
      17'd50663: data = 8'h00;
      17'd50664: data = 8'h00;
      17'd50665: data = 8'h01;
      17'd50666: data = 8'h01;
      17'd50667: data = 8'h01;
      17'd50668: data = 8'h00;
      17'd50669: data = 8'hfe;
      17'd50670: data = 8'hfe;
      17'd50671: data = 8'hfe;
      17'd50672: data = 8'hfd;
      17'd50673: data = 8'hfd;
      17'd50674: data = 8'hfd;
      17'd50675: data = 8'hfe;
      17'd50676: data = 8'hfe;
      17'd50677: data = 8'hfe;
      17'd50678: data = 8'hfe;
      17'd50679: data = 8'h00;
      17'd50680: data = 8'h00;
      17'd50681: data = 8'h00;
      17'd50682: data = 8'h00;
      17'd50683: data = 8'h01;
      17'd50684: data = 8'h00;
      17'd50685: data = 8'h00;
      17'd50686: data = 8'h00;
      17'd50687: data = 8'hfe;
      17'd50688: data = 8'hfd;
      17'd50689: data = 8'hfe;
      17'd50690: data = 8'h00;
      17'd50691: data = 8'hfe;
      17'd50692: data = 8'hfd;
      17'd50693: data = 8'hfe;
      17'd50694: data = 8'h00;
      17'd50695: data = 8'h00;
      17'd50696: data = 8'h00;
      17'd50697: data = 8'h00;
      17'd50698: data = 8'h01;
      17'd50699: data = 8'h01;
      17'd50700: data = 8'h00;
      17'd50701: data = 8'h00;
      17'd50702: data = 8'hfe;
      17'd50703: data = 8'hfd;
      17'd50704: data = 8'hfd;
      17'd50705: data = 8'hfd;
      17'd50706: data = 8'hfe;
      17'd50707: data = 8'hfe;
      17'd50708: data = 8'hfd;
      17'd50709: data = 8'hfe;
      17'd50710: data = 8'h00;
      17'd50711: data = 8'h00;
      17'd50712: data = 8'h00;
      17'd50713: data = 8'h01;
      17'd50714: data = 8'h01;
      17'd50715: data = 8'hfe;
      17'd50716: data = 8'h00;
      17'd50717: data = 8'h00;
      17'd50718: data = 8'hfd;
      17'd50719: data = 8'hfd;
      17'd50720: data = 8'hfd;
      17'd50721: data = 8'hfd;
      17'd50722: data = 8'hfd;
      17'd50723: data = 8'hfd;
      17'd50724: data = 8'hfd;
      17'd50725: data = 8'hfe;
      17'd50726: data = 8'h00;
      17'd50727: data = 8'h00;
      17'd50728: data = 8'h01;
      17'd50729: data = 8'h01;
      17'd50730: data = 8'h00;
      17'd50731: data = 8'h00;
      17'd50732: data = 8'h00;
      17'd50733: data = 8'hfe;
      17'd50734: data = 8'hfd;
      17'd50735: data = 8'hfe;
      17'd50736: data = 8'hfe;
      17'd50737: data = 8'hfd;
      17'd50738: data = 8'hfd;
      17'd50739: data = 8'hfd;
      17'd50740: data = 8'hfd;
      17'd50741: data = 8'hfe;
      17'd50742: data = 8'hfe;
      17'd50743: data = 8'h00;
      17'd50744: data = 8'hfe;
      17'd50745: data = 8'hfe;
      17'd50746: data = 8'hfe;
      17'd50747: data = 8'h00;
      17'd50748: data = 8'h00;
      17'd50749: data = 8'hfe;
      17'd50750: data = 8'hfe;
      17'd50751: data = 8'hfe;
      17'd50752: data = 8'hfe;
      17'd50753: data = 8'hfe;
      17'd50754: data = 8'hfd;
      17'd50755: data = 8'hfd;
      17'd50756: data = 8'hfe;
      17'd50757: data = 8'h00;
      17'd50758: data = 8'hfe;
      17'd50759: data = 8'h00;
      17'd50760: data = 8'h00;
      17'd50761: data = 8'h01;
      17'd50762: data = 8'h02;
      17'd50763: data = 8'h01;
      17'd50764: data = 8'h01;
      17'd50765: data = 8'h00;
      17'd50766: data = 8'hfe;
      17'd50767: data = 8'hfe;
      17'd50768: data = 8'hfd;
      17'd50769: data = 8'hfd;
      17'd50770: data = 8'hfd;
      17'd50771: data = 8'hfd;
      17'd50772: data = 8'hfd;
      17'd50773: data = 8'hfe;
      17'd50774: data = 8'hfe;
      17'd50775: data = 8'hfe;
      17'd50776: data = 8'h00;
      17'd50777: data = 8'h00;
      17'd50778: data = 8'h00;
      17'd50779: data = 8'h00;
      17'd50780: data = 8'h00;
      17'd50781: data = 8'h00;
      17'd50782: data = 8'hfe;
      17'd50783: data = 8'hfd;
      17'd50784: data = 8'hfd;
      17'd50785: data = 8'hfe;
      17'd50786: data = 8'hfd;
      17'd50787: data = 8'hfe;
      17'd50788: data = 8'hfe;
      17'd50789: data = 8'h00;
      17'd50790: data = 8'h00;
      17'd50791: data = 8'h00;
      17'd50792: data = 8'h01;
      17'd50793: data = 8'h01;
      17'd50794: data = 8'h00;
      17'd50795: data = 8'h00;
      17'd50796: data = 8'h01;
      17'd50797: data = 8'h01;
      17'd50798: data = 8'h00;
      17'd50799: data = 8'h00;
      17'd50800: data = 8'h00;
      17'd50801: data = 8'h00;
      17'd50802: data = 8'h00;
      17'd50803: data = 8'h00;
      17'd50804: data = 8'h00;
      17'd50805: data = 8'h00;
      17'd50806: data = 8'h00;
      17'd50807: data = 8'h01;
      17'd50808: data = 8'h01;
      17'd50809: data = 8'h01;
      17'd50810: data = 8'h02;
      17'd50811: data = 8'h02;
      17'd50812: data = 8'h02;
      17'd50813: data = 8'h02;
      17'd50814: data = 8'h01;
      17'd50815: data = 8'h01;
      17'd50816: data = 8'h00;
      17'd50817: data = 8'hfe;
      17'd50818: data = 8'h00;
      17'd50819: data = 8'hfe;
      17'd50820: data = 8'hfe;
      17'd50821: data = 8'h00;
      17'd50822: data = 8'h00;
      17'd50823: data = 8'h01;
      17'd50824: data = 8'hfe;
      17'd50825: data = 8'h00;
      17'd50826: data = 8'h01;
      17'd50827: data = 8'h00;
      17'd50828: data = 8'h00;
      17'd50829: data = 8'h00;
      17'd50830: data = 8'h01;
      17'd50831: data = 8'h00;
      17'd50832: data = 8'h00;
      17'd50833: data = 8'hfd;
      17'd50834: data = 8'hfd;
      17'd50835: data = 8'h00;
      17'd50836: data = 8'hfd;
      17'd50837: data = 8'hfe;
      17'd50838: data = 8'h00;
      17'd50839: data = 8'h00;
      17'd50840: data = 8'h00;
      17'd50841: data = 8'h01;
      17'd50842: data = 8'h01;
      17'd50843: data = 8'h01;
      17'd50844: data = 8'hfe;
      17'd50845: data = 8'hfe;
      17'd50846: data = 8'h00;
      17'd50847: data = 8'h00;
      17'd50848: data = 8'hfd;
      17'd50849: data = 8'hfd;
      17'd50850: data = 8'hfe;
      17'd50851: data = 8'hfd;
      17'd50852: data = 8'hfd;
      17'd50853: data = 8'hfc;
      17'd50854: data = 8'hfc;
      17'd50855: data = 8'hfe;
      17'd50856: data = 8'hfe;
      17'd50857: data = 8'hfe;
      17'd50858: data = 8'h00;
      17'd50859: data = 8'h00;
      17'd50860: data = 8'h00;
      17'd50861: data = 8'h00;
      17'd50862: data = 8'h00;
      17'd50863: data = 8'hfe;
      17'd50864: data = 8'hfd;
      17'd50865: data = 8'hfc;
      17'd50866: data = 8'hfc;
      17'd50867: data = 8'hfd;
      17'd50868: data = 8'hfc;
      17'd50869: data = 8'hfc;
      17'd50870: data = 8'hfe;
      17'd50871: data = 8'hfe;
      17'd50872: data = 8'hfe;
      17'd50873: data = 8'h00;
      17'd50874: data = 8'h01;
      17'd50875: data = 8'h01;
      17'd50876: data = 8'h00;
      17'd50877: data = 8'hfe;
      17'd50878: data = 8'hfd;
      17'd50879: data = 8'hfd;
      17'd50880: data = 8'hfd;
      17'd50881: data = 8'hfc;
      17'd50882: data = 8'hfd;
      17'd50883: data = 8'hfd;
      17'd50884: data = 8'hfc;
      17'd50885: data = 8'hfe;
      17'd50886: data = 8'h00;
      17'd50887: data = 8'hfe;
      17'd50888: data = 8'h00;
      17'd50889: data = 8'h00;
      17'd50890: data = 8'h00;
      17'd50891: data = 8'h00;
      17'd50892: data = 8'h00;
      17'd50893: data = 8'hfe;
      17'd50894: data = 8'hfd;
      17'd50895: data = 8'hfd;
      17'd50896: data = 8'hfd;
      17'd50897: data = 8'hfc;
      17'd50898: data = 8'hfc;
      17'd50899: data = 8'hfc;
      17'd50900: data = 8'hfd;
      17'd50901: data = 8'hfe;
      17'd50902: data = 8'hfe;
      17'd50903: data = 8'hfe;
      17'd50904: data = 8'h00;
      17'd50905: data = 8'h01;
      17'd50906: data = 8'h00;
      17'd50907: data = 8'h01;
      17'd50908: data = 8'h00;
      17'd50909: data = 8'hfe;
      17'd50910: data = 8'hfe;
      17'd50911: data = 8'hfd;
      17'd50912: data = 8'hfd;
      17'd50913: data = 8'hfd;
      17'd50914: data = 8'hfd;
      17'd50915: data = 8'hfe;
      17'd50916: data = 8'hfe;
      17'd50917: data = 8'hfe;
      17'd50918: data = 8'h00;
      17'd50919: data = 8'h00;
      17'd50920: data = 8'h00;
      17'd50921: data = 8'h00;
      17'd50922: data = 8'hfe;
      17'd50923: data = 8'hfd;
      17'd50924: data = 8'hfd;
      17'd50925: data = 8'hfd;
      17'd50926: data = 8'hfd;
      17'd50927: data = 8'hfe;
      17'd50928: data = 8'hfe;
      17'd50929: data = 8'hfe;
      17'd50930: data = 8'h00;
      17'd50931: data = 8'h00;
      17'd50932: data = 8'h00;
      17'd50933: data = 8'h00;
      17'd50934: data = 8'h00;
      17'd50935: data = 8'hfe;
      17'd50936: data = 8'hfd;
      17'd50937: data = 8'hfe;
      17'd50938: data = 8'hfe;
      17'd50939: data = 8'h00;
      17'd50940: data = 8'hfe;
      17'd50941: data = 8'hfe;
      17'd50942: data = 8'h00;
      17'd50943: data = 8'h00;
      17'd50944: data = 8'h02;
      17'd50945: data = 8'h01;
      17'd50946: data = 8'h01;
      17'd50947: data = 8'h01;
      17'd50948: data = 8'h01;
      17'd50949: data = 8'h00;
      17'd50950: data = 8'hfe;
      17'd50951: data = 8'h00;
      17'd50952: data = 8'hfe;
      17'd50953: data = 8'hfe;
      17'd50954: data = 8'hfd;
      17'd50955: data = 8'hfe;
      17'd50956: data = 8'hfe;
      17'd50957: data = 8'h00;
      17'd50958: data = 8'h01;
      17'd50959: data = 8'h01;
      17'd50960: data = 8'h01;
      17'd50961: data = 8'h01;
      17'd50962: data = 8'h00;
      17'd50963: data = 8'h00;
      17'd50964: data = 8'h00;
      17'd50965: data = 8'hfe;
      17'd50966: data = 8'hfe;
      17'd50967: data = 8'hfd;
      17'd50968: data = 8'hfe;
      17'd50969: data = 8'hfe;
      17'd50970: data = 8'h00;
      17'd50971: data = 8'h00;
      17'd50972: data = 8'h01;
      17'd50973: data = 8'h02;
      17'd50974: data = 8'h01;
      17'd50975: data = 8'h01;
      17'd50976: data = 8'h00;
      17'd50977: data = 8'h00;
      17'd50978: data = 8'h00;
      17'd50979: data = 8'hfe;
      17'd50980: data = 8'hfd;
      17'd50981: data = 8'hfd;
      17'd50982: data = 8'hfe;
      17'd50983: data = 8'hfe;
      17'd50984: data = 8'hfe;
      17'd50985: data = 8'hfd;
      17'd50986: data = 8'hfe;
      17'd50987: data = 8'hfe;
      17'd50988: data = 8'h00;
      17'd50989: data = 8'h00;
      17'd50990: data = 8'h00;
      17'd50991: data = 8'h00;
      17'd50992: data = 8'h00;
      17'd50993: data = 8'hfe;
      17'd50994: data = 8'hfe;
      17'd50995: data = 8'hfe;
      17'd50996: data = 8'hfe;
      17'd50997: data = 8'hfe;
      17'd50998: data = 8'hfe;
      17'd50999: data = 8'h00;
      17'd51000: data = 8'h00;
      17'd51001: data = 8'h01;
      17'd51002: data = 8'h01;
      17'd51003: data = 8'h01;
      17'd51004: data = 8'h01;
      17'd51005: data = 8'h01;
      17'd51006: data = 8'h00;
      17'd51007: data = 8'hfe;
      17'd51008: data = 8'h00;
      17'd51009: data = 8'hfe;
      17'd51010: data = 8'hfe;
      17'd51011: data = 8'hfe;
      17'd51012: data = 8'h00;
      17'd51013: data = 8'h01;
      17'd51014: data = 8'hfe;
      17'd51015: data = 8'h00;
      17'd51016: data = 8'h01;
      17'd51017: data = 8'h01;
      17'd51018: data = 8'h01;
      17'd51019: data = 8'h00;
      17'd51020: data = 8'h01;
      17'd51021: data = 8'h01;
      17'd51022: data = 8'h00;
      17'd51023: data = 8'h00;
      17'd51024: data = 8'h00;
      17'd51025: data = 8'h00;
      17'd51026: data = 8'hfd;
      17'd51027: data = 8'hfd;
      17'd51028: data = 8'hfe;
      17'd51029: data = 8'h00;
      17'd51030: data = 8'hfe;
      17'd51031: data = 8'h00;
      17'd51032: data = 8'h00;
      17'd51033: data = 8'h01;
      17'd51034: data = 8'h01;
      17'd51035: data = 8'hfe;
      17'd51036: data = 8'hfd;
      17'd51037: data = 8'hfe;
      17'd51038: data = 8'hfe;
      17'd51039: data = 8'hfd;
      17'd51040: data = 8'h00;
      17'd51041: data = 8'h00;
      17'd51042: data = 8'h00;
      17'd51043: data = 8'h01;
      17'd51044: data = 8'h00;
      17'd51045: data = 8'h01;
      17'd51046: data = 8'h00;
      17'd51047: data = 8'hfe;
      17'd51048: data = 8'h00;
      17'd51049: data = 8'h00;
      17'd51050: data = 8'h00;
      17'd51051: data = 8'h00;
      17'd51052: data = 8'h00;
      17'd51053: data = 8'hfe;
      17'd51054: data = 8'hfd;
      17'd51055: data = 8'hfd;
      17'd51056: data = 8'hfe;
      17'd51057: data = 8'hfe;
      17'd51058: data = 8'hfe;
      17'd51059: data = 8'h01;
      17'd51060: data = 8'h02;
      17'd51061: data = 8'h02;
      17'd51062: data = 8'h02;
      17'd51063: data = 8'h00;
      17'd51064: data = 8'h00;
      17'd51065: data = 8'h00;
      17'd51066: data = 8'hfd;
      17'd51067: data = 8'hfd;
      17'd51068: data = 8'hfd;
      17'd51069: data = 8'hfd;
      17'd51070: data = 8'hfe;
      17'd51071: data = 8'hfe;
      17'd51072: data = 8'hfe;
      17'd51073: data = 8'h00;
      17'd51074: data = 8'h00;
      17'd51075: data = 8'h00;
      17'd51076: data = 8'h01;
      17'd51077: data = 8'h01;
      17'd51078: data = 8'h00;
      17'd51079: data = 8'h00;
      17'd51080: data = 8'hfe;
      17'd51081: data = 8'hfd;
      17'd51082: data = 8'hfd;
      17'd51083: data = 8'hfd;
      17'd51084: data = 8'hfe;
      17'd51085: data = 8'hfe;
      17'd51086: data = 8'h00;
      17'd51087: data = 8'h00;
      17'd51088: data = 8'h00;
      17'd51089: data = 8'h01;
      17'd51090: data = 8'h01;
      17'd51091: data = 8'h00;
      17'd51092: data = 8'h00;
      17'd51093: data = 8'hfe;
      17'd51094: data = 8'hfe;
      17'd51095: data = 8'hfe;
      17'd51096: data = 8'hfd;
      17'd51097: data = 8'h00;
      17'd51098: data = 8'hfe;
      17'd51099: data = 8'hfe;
      17'd51100: data = 8'h01;
      17'd51101: data = 8'h01;
      17'd51102: data = 8'h01;
      17'd51103: data = 8'h01;
      17'd51104: data = 8'h01;
      17'd51105: data = 8'h01;
      17'd51106: data = 8'h01;
      17'd51107: data = 8'h00;
      17'd51108: data = 8'hfe;
      17'd51109: data = 8'hfe;
      17'd51110: data = 8'hfe;
      17'd51111: data = 8'hfd;
      17'd51112: data = 8'hfd;
      17'd51113: data = 8'hfd;
      17'd51114: data = 8'hfd;
      17'd51115: data = 8'hfe;
      17'd51116: data = 8'h01;
      17'd51117: data = 8'h01;
      17'd51118: data = 8'h00;
      17'd51119: data = 8'h02;
      17'd51120: data = 8'h01;
      17'd51121: data = 8'h00;
      17'd51122: data = 8'h00;
      17'd51123: data = 8'hfe;
      17'd51124: data = 8'hfe;
      17'd51125: data = 8'hfe;
      17'd51126: data = 8'h00;
      17'd51127: data = 8'hfe;
      17'd51128: data = 8'hfe;
      17'd51129: data = 8'h00;
      17'd51130: data = 8'h01;
      17'd51131: data = 8'h00;
      17'd51132: data = 8'h01;
      17'd51133: data = 8'h01;
      17'd51134: data = 8'h01;
      17'd51135: data = 8'h01;
      17'd51136: data = 8'h00;
      17'd51137: data = 8'hfe;
      17'd51138: data = 8'hfe;
      17'd51139: data = 8'hfe;
      17'd51140: data = 8'hfd;
      17'd51141: data = 8'hfd;
      17'd51142: data = 8'hfd;
      17'd51143: data = 8'hfe;
      17'd51144: data = 8'hfd;
      17'd51145: data = 8'hfe;
      17'd51146: data = 8'h00;
      17'd51147: data = 8'hfe;
      17'd51148: data = 8'h00;
      17'd51149: data = 8'h01;
      17'd51150: data = 8'h00;
      17'd51151: data = 8'hfe;
      17'd51152: data = 8'hfe;
      17'd51153: data = 8'h00;
      17'd51154: data = 8'hfe;
      17'd51155: data = 8'hfd;
      17'd51156: data = 8'hfd;
      17'd51157: data = 8'hfd;
      17'd51158: data = 8'hfd;
      17'd51159: data = 8'hfe;
      17'd51160: data = 8'hfe;
      17'd51161: data = 8'hfe;
      17'd51162: data = 8'h00;
      17'd51163: data = 8'h01;
      17'd51164: data = 8'h01;
      17'd51165: data = 8'h01;
      17'd51166: data = 8'h01;
      17'd51167: data = 8'hfe;
      17'd51168: data = 8'hfe;
      17'd51169: data = 8'hfe;
      17'd51170: data = 8'hfe;
      17'd51171: data = 8'hfd;
      17'd51172: data = 8'hfd;
      17'd51173: data = 8'hfe;
      17'd51174: data = 8'hfe;
      17'd51175: data = 8'h00;
      17'd51176: data = 8'h00;
      17'd51177: data = 8'h00;
      17'd51178: data = 8'h01;
      17'd51179: data = 8'h00;
      17'd51180: data = 8'h00;
      17'd51181: data = 8'hfe;
      17'd51182: data = 8'hfe;
      17'd51183: data = 8'hfe;
      17'd51184: data = 8'hfd;
      17'd51185: data = 8'hfd;
      17'd51186: data = 8'hfd;
      17'd51187: data = 8'hfd;
      17'd51188: data = 8'hfd;
      17'd51189: data = 8'h00;
      17'd51190: data = 8'h01;
      17'd51191: data = 8'h01;
      17'd51192: data = 8'h02;
      17'd51193: data = 8'h02;
      17'd51194: data = 8'h01;
      17'd51195: data = 8'h01;
      17'd51196: data = 8'hfe;
      17'd51197: data = 8'hfd;
      17'd51198: data = 8'hfd;
      17'd51199: data = 8'hfd;
      17'd51200: data = 8'hfc;
      17'd51201: data = 8'hfc;
      17'd51202: data = 8'hfe;
      17'd51203: data = 8'hfe;
      17'd51204: data = 8'h00;
      17'd51205: data = 8'h01;
      17'd51206: data = 8'h01;
      17'd51207: data = 8'h01;
      17'd51208: data = 8'h01;
      17'd51209: data = 8'h00;
      17'd51210: data = 8'hfe;
      17'd51211: data = 8'hfe;
      17'd51212: data = 8'hfd;
      17'd51213: data = 8'hfc;
      17'd51214: data = 8'hfd;
      17'd51215: data = 8'hfc;
      17'd51216: data = 8'hfd;
      17'd51217: data = 8'hfe;
      17'd51218: data = 8'hfd;
      17'd51219: data = 8'h00;
      17'd51220: data = 8'h01;
      17'd51221: data = 8'h01;
      17'd51222: data = 8'h01;
      17'd51223: data = 8'h01;
      17'd51224: data = 8'h01;
      17'd51225: data = 8'hfe;
      17'd51226: data = 8'h00;
      17'd51227: data = 8'h00;
      17'd51228: data = 8'hfd;
      17'd51229: data = 8'hfd;
      17'd51230: data = 8'hfd;
      17'd51231: data = 8'hfd;
      17'd51232: data = 8'h00;
      17'd51233: data = 8'h01;
      17'd51234: data = 8'hfe;
      17'd51235: data = 8'h01;
      17'd51236: data = 8'h04;
      17'd51237: data = 8'h02;
      17'd51238: data = 8'h01;
      17'd51239: data = 8'h00;
      17'd51240: data = 8'h00;
      17'd51241: data = 8'hfe;
      17'd51242: data = 8'hfe;
      17'd51243: data = 8'hfd;
      17'd51244: data = 8'hfd;
      17'd51245: data = 8'hfd;
      17'd51246: data = 8'hfe;
      17'd51247: data = 8'hfe;
      17'd51248: data = 8'h00;
      17'd51249: data = 8'h01;
      17'd51250: data = 8'h00;
      17'd51251: data = 8'h02;
      17'd51252: data = 8'h04;
      17'd51253: data = 8'h02;
      17'd51254: data = 8'h01;
      17'd51255: data = 8'h00;
      17'd51256: data = 8'h00;
      17'd51257: data = 8'hfe;
      17'd51258: data = 8'hfe;
      17'd51259: data = 8'hfd;
      17'd51260: data = 8'hfd;
      17'd51261: data = 8'hfe;
      17'd51262: data = 8'h00;
      17'd51263: data = 8'h02;
      17'd51264: data = 8'h04;
      17'd51265: data = 8'h04;
      17'd51266: data = 8'h04;
      17'd51267: data = 8'h02;
      17'd51268: data = 8'h01;
      17'd51269: data = 8'h01;
      17'd51270: data = 8'h00;
      17'd51271: data = 8'hfd;
      17'd51272: data = 8'hfd;
      17'd51273: data = 8'hfd;
      17'd51274: data = 8'hfe;
      17'd51275: data = 8'hfe;
      17'd51276: data = 8'hfe;
      17'd51277: data = 8'h00;
      17'd51278: data = 8'h02;
      17'd51279: data = 8'h02;
      17'd51280: data = 8'h01;
      17'd51281: data = 8'h02;
      17'd51282: data = 8'h01;
      17'd51283: data = 8'h01;
      17'd51284: data = 8'hfe;
      17'd51285: data = 8'hfd;
      17'd51286: data = 8'hfc;
      17'd51287: data = 8'hfc;
      17'd51288: data = 8'hfc;
      17'd51289: data = 8'hfc;
      17'd51290: data = 8'hfd;
      17'd51291: data = 8'hfe;
      17'd51292: data = 8'h00;
      17'd51293: data = 8'h01;
      17'd51294: data = 8'h01;
      17'd51295: data = 8'h02;
      17'd51296: data = 8'h02;
      17'd51297: data = 8'h01;
      17'd51298: data = 8'h00;
      17'd51299: data = 8'hfe;
      17'd51300: data = 8'hfd;
      17'd51301: data = 8'hfd;
      17'd51302: data = 8'hfd;
      17'd51303: data = 8'hfc;
      17'd51304: data = 8'hfd;
      17'd51305: data = 8'hfe;
      17'd51306: data = 8'h01;
      17'd51307: data = 8'h01;
      17'd51308: data = 8'h01;
      17'd51309: data = 8'h01;
      17'd51310: data = 8'h01;
      17'd51311: data = 8'h01;
      17'd51312: data = 8'h00;
      17'd51313: data = 8'h01;
      17'd51314: data = 8'h00;
      17'd51315: data = 8'hfe;
      17'd51316: data = 8'hfe;
      17'd51317: data = 8'hfe;
      17'd51318: data = 8'hfd;
      17'd51319: data = 8'hfe;
      17'd51320: data = 8'h00;
      17'd51321: data = 8'h00;
      17'd51322: data = 8'h00;
      17'd51323: data = 8'h01;
      17'd51324: data = 8'h00;
      17'd51325: data = 8'h01;
      17'd51326: data = 8'h00;
      17'd51327: data = 8'h00;
      17'd51328: data = 8'hfe;
      17'd51329: data = 8'hfd;
      17'd51330: data = 8'hfe;
      17'd51331: data = 8'hfd;
      17'd51332: data = 8'hfd;
      17'd51333: data = 8'hfe;
      17'd51334: data = 8'hfe;
      17'd51335: data = 8'hfe;
      17'd51336: data = 8'h00;
      17'd51337: data = 8'h01;
      17'd51338: data = 8'h01;
      17'd51339: data = 8'h01;
      17'd51340: data = 8'h01;
      17'd51341: data = 8'h01;
      17'd51342: data = 8'h00;
      17'd51343: data = 8'hfe;
      17'd51344: data = 8'hfe;
      17'd51345: data = 8'hfd;
      17'd51346: data = 8'hfd;
      17'd51347: data = 8'hfe;
      17'd51348: data = 8'hfe;
      17'd51349: data = 8'h00;
      17'd51350: data = 8'h01;
      17'd51351: data = 8'h01;
      17'd51352: data = 8'h01;
      17'd51353: data = 8'h02;
      17'd51354: data = 8'h01;
      17'd51355: data = 8'h02;
      17'd51356: data = 8'h01;
      17'd51357: data = 8'h00;
      17'd51358: data = 8'h00;
      17'd51359: data = 8'hfd;
      17'd51360: data = 8'hfd;
      17'd51361: data = 8'hfe;
      17'd51362: data = 8'hfd;
      17'd51363: data = 8'hfd;
      17'd51364: data = 8'hfe;
      17'd51365: data = 8'h01;
      17'd51366: data = 8'h01;
      17'd51367: data = 8'h01;
      17'd51368: data = 8'h02;
      17'd51369: data = 8'h00;
      17'd51370: data = 8'h00;
      17'd51371: data = 8'h00;
      17'd51372: data = 8'hfe;
      17'd51373: data = 8'hfe;
      17'd51374: data = 8'hfe;
      17'd51375: data = 8'hfe;
      17'd51376: data = 8'hfe;
      17'd51377: data = 8'hfe;
      17'd51378: data = 8'h01;
      17'd51379: data = 8'h00;
      17'd51380: data = 8'hfe;
      17'd51381: data = 8'h00;
      17'd51382: data = 8'hfe;
      17'd51383: data = 8'h00;
      17'd51384: data = 8'hfe;
      17'd51385: data = 8'hfe;
      17'd51386: data = 8'hfe;
      17'd51387: data = 8'hfe;
      17'd51388: data = 8'hfe;
      17'd51389: data = 8'hfe;
      17'd51390: data = 8'h00;
      17'd51391: data = 8'hfe;
      17'd51392: data = 8'h00;
      17'd51393: data = 8'h00;
      17'd51394: data = 8'hfe;
      17'd51395: data = 8'h00;
      17'd51396: data = 8'hfe;
      17'd51397: data = 8'hfe;
      17'd51398: data = 8'hfe;
      17'd51399: data = 8'hfd;
      17'd51400: data = 8'hfd;
      17'd51401: data = 8'hfd;
      17'd51402: data = 8'hfe;
      17'd51403: data = 8'h01;
      17'd51404: data = 8'h00;
      17'd51405: data = 8'h00;
      17'd51406: data = 8'h01;
      17'd51407: data = 8'h01;
      17'd51408: data = 8'h01;
      17'd51409: data = 8'h00;
      17'd51410: data = 8'hfe;
      17'd51411: data = 8'h00;
      17'd51412: data = 8'hfe;
      17'd51413: data = 8'hfd;
      17'd51414: data = 8'hfe;
      17'd51415: data = 8'hfe;
      17'd51416: data = 8'hfe;
      17'd51417: data = 8'hfe;
      17'd51418: data = 8'hfe;
      17'd51419: data = 8'h00;
      17'd51420: data = 8'h01;
      17'd51421: data = 8'h01;
      17'd51422: data = 8'h00;
      17'd51423: data = 8'h01;
      17'd51424: data = 8'h01;
      17'd51425: data = 8'hfe;
      17'd51426: data = 8'hfd;
      17'd51427: data = 8'hfe;
      17'd51428: data = 8'hfd;
      17'd51429: data = 8'hfd;
      17'd51430: data = 8'hfd;
      17'd51431: data = 8'hfd;
      17'd51432: data = 8'hfd;
      17'd51433: data = 8'hfe;
      17'd51434: data = 8'hfe;
      17'd51435: data = 8'h00;
      17'd51436: data = 8'h00;
      17'd51437: data = 8'h00;
      17'd51438: data = 8'h00;
      17'd51439: data = 8'h00;
      17'd51440: data = 8'h00;
      17'd51441: data = 8'hfe;
      17'd51442: data = 8'hfe;
      17'd51443: data = 8'hfe;
      17'd51444: data = 8'hfe;
      17'd51445: data = 8'hfd;
      17'd51446: data = 8'hfe;
      17'd51447: data = 8'hfe;
      17'd51448: data = 8'h00;
      17'd51449: data = 8'hfe;
      17'd51450: data = 8'hfe;
      17'd51451: data = 8'h00;
      17'd51452: data = 8'hfe;
      17'd51453: data = 8'h00;
      17'd51454: data = 8'hfe;
      17'd51455: data = 8'h00;
      17'd51456: data = 8'h00;
      17'd51457: data = 8'h00;
      17'd51458: data = 8'hfe;
      17'd51459: data = 8'hfe;
      17'd51460: data = 8'hfe;
      17'd51461: data = 8'hfd;
      17'd51462: data = 8'hfe;
      17'd51463: data = 8'h00;
      17'd51464: data = 8'h00;
      17'd51465: data = 8'h00;
      17'd51466: data = 8'h01;
      17'd51467: data = 8'h01;
      17'd51468: data = 8'h01;
      17'd51469: data = 8'h01;
      17'd51470: data = 8'h00;
      17'd51471: data = 8'hfe;
      17'd51472: data = 8'h00;
      17'd51473: data = 8'h00;
      17'd51474: data = 8'hfe;
      17'd51475: data = 8'hfe;
      17'd51476: data = 8'h00;
      17'd51477: data = 8'hfe;
      17'd51478: data = 8'hfe;
      17'd51479: data = 8'hfe;
      17'd51480: data = 8'h01;
      17'd51481: data = 8'h01;
      17'd51482: data = 8'h01;
      17'd51483: data = 8'h04;
      17'd51484: data = 8'h02;
      17'd51485: data = 8'h02;
      17'd51486: data = 8'h01;
      17'd51487: data = 8'h00;
      17'd51488: data = 8'h00;
      17'd51489: data = 8'hfe;
      17'd51490: data = 8'hfe;
      17'd51491: data = 8'hfe;
      17'd51492: data = 8'hfe;
      17'd51493: data = 8'h00;
      17'd51494: data = 8'h01;
      17'd51495: data = 8'h00;
      17'd51496: data = 8'h01;
      17'd51497: data = 8'h01;
      17'd51498: data = 8'h02;
      17'd51499: data = 8'h01;
      17'd51500: data = 8'h00;
      17'd51501: data = 8'hfe;
      17'd51502: data = 8'hfd;
      17'd51503: data = 8'hfe;
      17'd51504: data = 8'hfd;
      17'd51505: data = 8'hfe;
      17'd51506: data = 8'h00;
      17'd51507: data = 8'h01;
      17'd51508: data = 8'h02;
      17'd51509: data = 8'h01;
      17'd51510: data = 8'h01;
      17'd51511: data = 8'h01;
      17'd51512: data = 8'h01;
      17'd51513: data = 8'h00;
      17'd51514: data = 8'h02;
      17'd51515: data = 8'h01;
      17'd51516: data = 8'h00;
      17'd51517: data = 8'h01;
      17'd51518: data = 8'h00;
      17'd51519: data = 8'hfe;
      17'd51520: data = 8'hfe;
      17'd51521: data = 8'hfe;
      17'd51522: data = 8'h01;
      17'd51523: data = 8'h00;
      17'd51524: data = 8'h00;
      17'd51525: data = 8'h01;
      17'd51526: data = 8'h01;
      17'd51527: data = 8'h01;
      17'd51528: data = 8'h00;
      17'd51529: data = 8'hfe;
      17'd51530: data = 8'h00;
      17'd51531: data = 8'h00;
      17'd51532: data = 8'hfe;
      17'd51533: data = 8'h00;
      17'd51534: data = 8'hfe;
      17'd51535: data = 8'h00;
      17'd51536: data = 8'h01;
      17'd51537: data = 8'h00;
      17'd51538: data = 8'h00;
      17'd51539: data = 8'h00;
      17'd51540: data = 8'h00;
      17'd51541: data = 8'h00;
      17'd51542: data = 8'h01;
      17'd51543: data = 8'h01;
      17'd51544: data = 8'h00;
      17'd51545: data = 8'h01;
      17'd51546: data = 8'h00;
      17'd51547: data = 8'h00;
      17'd51548: data = 8'h00;
      17'd51549: data = 8'h00;
      17'd51550: data = 8'h00;
      17'd51551: data = 8'h00;
      17'd51552: data = 8'h01;
      17'd51553: data = 8'h01;
      17'd51554: data = 8'h01;
      17'd51555: data = 8'h01;
      17'd51556: data = 8'h01;
      17'd51557: data = 8'h00;
      17'd51558: data = 8'h00;
      17'd51559: data = 8'h00;
      17'd51560: data = 8'hfe;
      17'd51561: data = 8'h00;
      17'd51562: data = 8'h01;
      17'd51563: data = 8'hfe;
      17'd51564: data = 8'hfd;
      17'd51565: data = 8'hfe;
      17'd51566: data = 8'h00;
      17'd51567: data = 8'h00;
      17'd51568: data = 8'h00;
      17'd51569: data = 8'hfe;
      17'd51570: data = 8'h00;
      17'd51571: data = 8'h00;
      17'd51572: data = 8'h00;
      17'd51573: data = 8'hfe;
      17'd51574: data = 8'h00;
      17'd51575: data = 8'h00;
      17'd51576: data = 8'hfe;
      17'd51577: data = 8'hfe;
      17'd51578: data = 8'hfe;
      17'd51579: data = 8'h00;
      17'd51580: data = 8'h00;
      17'd51581: data = 8'hfe;
      17'd51582: data = 8'hfd;
      17'd51583: data = 8'hfd;
      17'd51584: data = 8'hfd;
      17'd51585: data = 8'hfd;
      17'd51586: data = 8'hfc;
      17'd51587: data = 8'hfc;
      17'd51588: data = 8'hfa;
      17'd51589: data = 8'hfc;
      17'd51590: data = 8'hfe;
      17'd51591: data = 8'h02;
      17'd51592: data = 8'h02;
      17'd51593: data = 8'h01;
      17'd51594: data = 8'h02;
      17'd51595: data = 8'h00;
      17'd51596: data = 8'h00;
      17'd51597: data = 8'h04;
      17'd51598: data = 8'h06;
      17'd51599: data = 8'h05;
      17'd51600: data = 8'h09;
      17'd51601: data = 8'h0a;
      17'd51602: data = 8'h02;
      17'd51603: data = 8'hfe;
      17'd51604: data = 8'hfd;
      17'd51605: data = 8'hf9;
      17'd51606: data = 8'hf6;
      17'd51607: data = 8'hfd;
      17'd51608: data = 8'hfd;
      17'd51609: data = 8'hfa;
      17'd51610: data = 8'hfd;
      17'd51611: data = 8'hfd;
      17'd51612: data = 8'h00;
      17'd51613: data = 8'h01;
      17'd51614: data = 8'hfe;
      17'd51615: data = 8'hfe;
      17'd51616: data = 8'hfc;
      17'd51617: data = 8'hfd;
      17'd51618: data = 8'h00;
      17'd51619: data = 8'h02;
      17'd51620: data = 8'h01;
      17'd51621: data = 8'hfe;
      17'd51622: data = 8'hfc;
      17'd51623: data = 8'hfc;
      17'd51624: data = 8'hfa;
      17'd51625: data = 8'hfc;
      17'd51626: data = 8'hfd;
      17'd51627: data = 8'hfd;
      17'd51628: data = 8'hfe;
      17'd51629: data = 8'h01;
      17'd51630: data = 8'h01;
      17'd51631: data = 8'h02;
      17'd51632: data = 8'h02;
      17'd51633: data = 8'h01;
      17'd51634: data = 8'h00;
      17'd51635: data = 8'h00;
      17'd51636: data = 8'hfe;
      17'd51637: data = 8'h01;
      17'd51638: data = 8'h01;
      17'd51639: data = 8'h02;
      17'd51640: data = 8'h02;
      17'd51641: data = 8'h00;
      17'd51642: data = 8'h00;
      17'd51643: data = 8'hfe;
      17'd51644: data = 8'hfd;
      17'd51645: data = 8'hfd;
      17'd51646: data = 8'hfe;
      17'd51647: data = 8'h00;
      17'd51648: data = 8'h00;
      17'd51649: data = 8'h01;
      17'd51650: data = 8'h01;
      17'd51651: data = 8'h00;
      17'd51652: data = 8'h00;
      17'd51653: data = 8'hfe;
      17'd51654: data = 8'hfe;
      17'd51655: data = 8'h01;
      17'd51656: data = 8'h01;
      17'd51657: data = 8'h01;
      17'd51658: data = 8'hfe;
      17'd51659: data = 8'h02;
      17'd51660: data = 8'h04;
      17'd51661: data = 8'hfe;
      17'd51662: data = 8'h01;
      17'd51663: data = 8'hfe;
      17'd51664: data = 8'hfd;
      17'd51665: data = 8'h01;
      17'd51666: data = 8'h01;
      17'd51667: data = 8'h02;
      17'd51668: data = 8'h00;
      17'd51669: data = 8'hfe;
      17'd51670: data = 8'hfe;
      17'd51671: data = 8'hfe;
      17'd51672: data = 8'hfe;
      17'd51673: data = 8'hfe;
      17'd51674: data = 8'hfe;
      17'd51675: data = 8'hfd;
      17'd51676: data = 8'h00;
      17'd51677: data = 8'hfe;
      17'd51678: data = 8'h01;
      17'd51679: data = 8'h01;
      17'd51680: data = 8'hfe;
      17'd51681: data = 8'hfd;
      17'd51682: data = 8'hfc;
      17'd51683: data = 8'hfc;
      17'd51684: data = 8'hfd;
      17'd51685: data = 8'hfe;
      17'd51686: data = 8'hfd;
      17'd51687: data = 8'h00;
      17'd51688: data = 8'h01;
      17'd51689: data = 8'hfd;
      17'd51690: data = 8'h00;
      17'd51691: data = 8'h00;
      17'd51692: data = 8'h00;
      17'd51693: data = 8'h00;
      17'd51694: data = 8'hfd;
      17'd51695: data = 8'hfc;
      17'd51696: data = 8'hfa;
      17'd51697: data = 8'hfc;
      17'd51698: data = 8'h02;
      17'd51699: data = 8'h01;
      17'd51700: data = 8'hfe;
      17'd51701: data = 8'h01;
      17'd51702: data = 8'h00;
      17'd51703: data = 8'h02;
      17'd51704: data = 8'h02;
      17'd51705: data = 8'hfe;
      17'd51706: data = 8'hfd;
      17'd51707: data = 8'hfa;
      17'd51708: data = 8'hfa;
      17'd51709: data = 8'hfd;
      17'd51710: data = 8'hf6;
      17'd51711: data = 8'hf9;
      17'd51712: data = 8'hf6;
      17'd51713: data = 8'hf9;
      17'd51714: data = 8'h00;
      17'd51715: data = 8'h00;
      17'd51716: data = 8'h01;
      17'd51717: data = 8'h00;
      17'd51718: data = 8'hfd;
      17'd51719: data = 8'hfe;
      17'd51720: data = 8'h05;
      17'd51721: data = 8'h05;
      17'd51722: data = 8'h04;
      17'd51723: data = 8'h00;
      17'd51724: data = 8'hfa;
      17'd51725: data = 8'hf9;
      17'd51726: data = 8'hfa;
      17'd51727: data = 8'hfa;
      17'd51728: data = 8'hfe;
      17'd51729: data = 8'h02;
      17'd51730: data = 8'h02;
      17'd51731: data = 8'h00;
      17'd51732: data = 8'h01;
      17'd51733: data = 8'h05;
      17'd51734: data = 8'h05;
      17'd51735: data = 8'h09;
      17'd51736: data = 8'h0a;
      17'd51737: data = 8'h09;
      17'd51738: data = 8'h04;
      17'd51739: data = 8'hfe;
      17'd51740: data = 8'h00;
      17'd51741: data = 8'hfd;
      17'd51742: data = 8'h00;
      17'd51743: data = 8'hfa;
      17'd51744: data = 8'hf4;
      17'd51745: data = 8'hf1;
      17'd51746: data = 8'heb;
      17'd51747: data = 8'hf2;
      17'd51748: data = 8'hf5;
      17'd51749: data = 8'hf9;
      17'd51750: data = 8'hfd;
      17'd51751: data = 8'hf6;
      17'd51752: data = 8'hef;
      17'd51753: data = 8'hf4;
      17'd51754: data = 8'hf5;
      17'd51755: data = 8'hfe;
      17'd51756: data = 8'h0c;
      17'd51757: data = 8'h0e;
      17'd51758: data = 8'h13;
      17'd51759: data = 8'h15;
      17'd51760: data = 8'h16;
      17'd51761: data = 8'h1b;
      17'd51762: data = 8'h1e;
      17'd51763: data = 8'h1f;
      17'd51764: data = 8'h1e;
      17'd51765: data = 8'h15;
      17'd51766: data = 8'h02;
      17'd51767: data = 8'hf2;
      17'd51768: data = 8'he4;
      17'd51769: data = 8'hdb;
      17'd51770: data = 8'he0;
      17'd51771: data = 8'hec;
      17'd51772: data = 8'hfc;
      17'd51773: data = 8'h06;
      17'd51774: data = 8'h09;
      17'd51775: data = 8'h06;
      17'd51776: data = 8'h02;
      17'd51777: data = 8'h02;
      17'd51778: data = 8'h05;
      17'd51779: data = 8'h12;
      17'd51780: data = 8'h23;
      17'd51781: data = 8'h2b;
      17'd51782: data = 8'h29;
      17'd51783: data = 8'h1b;
      17'd51784: data = 8'h04;
      17'd51785: data = 8'hf1;
      17'd51786: data = 8'he3;
      17'd51787: data = 8'hda;
      17'd51788: data = 8'he0;
      17'd51789: data = 8'he3;
      17'd51790: data = 8'he5;
      17'd51791: data = 8'heb;
      17'd51792: data = 8'he9;
      17'd51793: data = 8'he2;
      17'd51794: data = 8'hdc;
      17'd51795: data = 8'hdc;
      17'd51796: data = 8'he3;
      17'd51797: data = 8'hf4;
      17'd51798: data = 8'h02;
      17'd51799: data = 8'h13;
      17'd51800: data = 8'h1e;
      17'd51801: data = 8'h1c;
      17'd51802: data = 8'h16;
      17'd51803: data = 8'h11;
      17'd51804: data = 8'h0a;
      17'd51805: data = 8'h05;
      17'd51806: data = 8'h06;
      17'd51807: data = 8'h05;
      17'd51808: data = 8'h04;
      17'd51809: data = 8'h02;
      17'd51810: data = 8'hfd;
      17'd51811: data = 8'hf6;
      17'd51812: data = 8'hef;
      17'd51813: data = 8'hed;
      17'd51814: data = 8'hef;
      17'd51815: data = 8'hf4;
      17'd51816: data = 8'hfa;
      17'd51817: data = 8'h02;
      17'd51818: data = 8'h0c;
      17'd51819: data = 8'h11;
      17'd51820: data = 8'h15;
      17'd51821: data = 8'h19;
      17'd51822: data = 8'h16;
      17'd51823: data = 8'h13;
      17'd51824: data = 8'h0e;
      17'd51825: data = 8'h0a;
      17'd51826: data = 8'h06;
      17'd51827: data = 8'h04;
      17'd51828: data = 8'h04;
      17'd51829: data = 8'hfe;
      17'd51830: data = 8'hf9;
      17'd51831: data = 8'hf4;
      17'd51832: data = 8'heb;
      17'd51833: data = 8'he3;
      17'd51834: data = 8'he3;
      17'd51835: data = 8'he7;
      17'd51836: data = 8'hed;
      17'd51837: data = 8'hf9;
      17'd51838: data = 8'h02;
      17'd51839: data = 8'h06;
      17'd51840: data = 8'h0d;
      17'd51841: data = 8'h13;
      17'd51842: data = 8'h15;
      17'd51843: data = 8'h16;
      17'd51844: data = 8'h1c;
      17'd51845: data = 8'h1e;
      17'd51846: data = 8'h1b;
      17'd51847: data = 8'h19;
      17'd51848: data = 8'h13;
      17'd51849: data = 8'h0d;
      17'd51850: data = 8'h05;
      17'd51851: data = 8'hfc;
      17'd51852: data = 8'hf4;
      17'd51853: data = 8'hef;
      17'd51854: data = 8'he9;
      17'd51855: data = 8'he7;
      17'd51856: data = 8'heb;
      17'd51857: data = 8'he7;
      17'd51858: data = 8'hec;
      17'd51859: data = 8'hf1;
      17'd51860: data = 8'hf2;
      17'd51861: data = 8'hf2;
      17'd51862: data = 8'hf5;
      17'd51863: data = 8'hf6;
      17'd51864: data = 8'hf6;
      17'd51865: data = 8'hfc;
      17'd51866: data = 8'h01;
      17'd51867: data = 8'h01;
      17'd51868: data = 8'hfe;
      17'd51869: data = 8'hfd;
      17'd51870: data = 8'hfc;
      17'd51871: data = 8'hf6;
      17'd51872: data = 8'hf5;
      17'd51873: data = 8'hfa;
      17'd51874: data = 8'hfa;
      17'd51875: data = 8'hf9;
      17'd51876: data = 8'hfe;
      17'd51877: data = 8'h02;
      17'd51878: data = 8'h02;
      17'd51879: data = 8'h02;
      17'd51880: data = 8'h04;
      17'd51881: data = 8'h04;
      17'd51882: data = 8'h04;
      17'd51883: data = 8'h02;
      17'd51884: data = 8'h02;
      17'd51885: data = 8'h01;
      17'd51886: data = 8'h00;
      17'd51887: data = 8'hfe;
      17'd51888: data = 8'hf9;
      17'd51889: data = 8'hf5;
      17'd51890: data = 8'hf1;
      17'd51891: data = 8'hed;
      17'd51892: data = 8'hef;
      17'd51893: data = 8'hed;
      17'd51894: data = 8'hf2;
      17'd51895: data = 8'hf5;
      17'd51896: data = 8'hf5;
      17'd51897: data = 8'hf9;
      17'd51898: data = 8'hfc;
      17'd51899: data = 8'h00;
      17'd51900: data = 8'h02;
      17'd51901: data = 8'h04;
      17'd51902: data = 8'h05;
      17'd51903: data = 8'h05;
      17'd51904: data = 8'h06;
      17'd51905: data = 8'h09;
      17'd51906: data = 8'h06;
      17'd51907: data = 8'h05;
      17'd51908: data = 8'h00;
      17'd51909: data = 8'hfd;
      17'd51910: data = 8'hfd;
      17'd51911: data = 8'hfa;
      17'd51912: data = 8'hfd;
      17'd51913: data = 8'hf9;
      17'd51914: data = 8'hf5;
      17'd51915: data = 8'hf5;
      17'd51916: data = 8'hf2;
      17'd51917: data = 8'hf6;
      17'd51918: data = 8'hf6;
      17'd51919: data = 8'hf9;
      17'd51920: data = 8'hfd;
      17'd51921: data = 8'hfd;
      17'd51922: data = 8'h00;
      17'd51923: data = 8'h00;
      17'd51924: data = 8'h00;
      17'd51925: data = 8'h02;
      17'd51926: data = 8'h01;
      17'd51927: data = 8'h06;
      17'd51928: data = 8'h06;
      17'd51929: data = 8'h02;
      17'd51930: data = 8'h04;
      17'd51931: data = 8'hfe;
      17'd51932: data = 8'hfd;
      17'd51933: data = 8'hfe;
      17'd51934: data = 8'h00;
      17'd51935: data = 8'h01;
      17'd51936: data = 8'h02;
      17'd51937: data = 8'h01;
      17'd51938: data = 8'h02;
      17'd51939: data = 8'h00;
      17'd51940: data = 8'hfe;
      17'd51941: data = 8'h00;
      17'd51942: data = 8'h02;
      17'd51943: data = 8'h05;
      17'd51944: data = 8'h09;
      17'd51945: data = 8'h0d;
      17'd51946: data = 8'h04;
      17'd51947: data = 8'h0c;
      17'd51948: data = 8'h0e;
      17'd51949: data = 8'h06;
      17'd51950: data = 8'h04;
      17'd51951: data = 8'hfd;
      17'd51952: data = 8'hf2;
      17'd51953: data = 8'hf6;
      17'd51954: data = 8'hfd;
      17'd51955: data = 8'h02;
      17'd51956: data = 8'h09;
      17'd51957: data = 8'hfd;
      17'd51958: data = 8'hf5;
      17'd51959: data = 8'hfa;
      17'd51960: data = 8'hfe;
      17'd51961: data = 8'h02;
      17'd51962: data = 8'h0d;
      17'd51963: data = 8'h05;
      17'd51964: data = 8'hfc;
      17'd51965: data = 8'hfe;
      17'd51966: data = 8'h05;
      17'd51967: data = 8'h04;
      17'd51968: data = 8'h05;
      17'd51969: data = 8'h01;
      17'd51970: data = 8'hf9;
      17'd51971: data = 8'hf6;
      17'd51972: data = 8'hfd;
      17'd51973: data = 8'hfd;
      17'd51974: data = 8'hf6;
      17'd51975: data = 8'hf5;
      17'd51976: data = 8'hf6;
      17'd51977: data = 8'hf9;
      17'd51978: data = 8'hfe;
      17'd51979: data = 8'h05;
      17'd51980: data = 8'h02;
      17'd51981: data = 8'h00;
      17'd51982: data = 8'h05;
      17'd51983: data = 8'h11;
      17'd51984: data = 8'h19;
      17'd51985: data = 8'h22;
      17'd51986: data = 8'h27;
      17'd51987: data = 8'h2b;
      17'd51988: data = 8'h2b;
      17'd51989: data = 8'h26;
      17'd51990: data = 8'h1c;
      17'd51991: data = 8'h16;
      17'd51992: data = 8'h0d;
      17'd51993: data = 8'h0d;
      17'd51994: data = 8'h16;
      17'd51995: data = 8'h1a;
      17'd51996: data = 8'h16;
      17'd51997: data = 8'h13;
      17'd51998: data = 8'h01;
      17'd51999: data = 8'heb;
      17'd52000: data = 8'he5;
      17'd52001: data = 8'he4;
      17'd52002: data = 8'he3;
      17'd52003: data = 8'heb;
      17'd52004: data = 8'hf4;
      17'd52005: data = 8'hf1;
      17'd52006: data = 8'hec;
      17'd52007: data = 8'he3;
      17'd52008: data = 8'hd8;
      17'd52009: data = 8'hd8;
      17'd52010: data = 8'hd6;
      17'd52011: data = 8'hda;
      17'd52012: data = 8'hde;
      17'd52013: data = 8'he0;
      17'd52014: data = 8'he4;
      17'd52015: data = 8'he7;
      17'd52016: data = 8'he4;
      17'd52017: data = 8'he4;
      17'd52018: data = 8'he3;
      17'd52019: data = 8'he5;
      17'd52020: data = 8'hf1;
      17'd52021: data = 8'hfc;
      17'd52022: data = 8'h06;
      17'd52023: data = 8'h0d;
      17'd52024: data = 8'h0d;
      17'd52025: data = 8'h11;
      17'd52026: data = 8'h12;
      17'd52027: data = 8'h12;
      17'd52028: data = 8'h12;
      17'd52029: data = 8'h16;
      17'd52030: data = 8'h15;
      17'd52031: data = 8'h15;
      17'd52032: data = 8'h1e;
      17'd52033: data = 8'h1f;
      17'd52034: data = 8'h1c;
      17'd52035: data = 8'h1f;
      17'd52036: data = 8'h1b;
      17'd52037: data = 8'h13;
      17'd52038: data = 8'h11;
      17'd52039: data = 8'h0e;
      17'd52040: data = 8'h0c;
      17'd52041: data = 8'h09;
      17'd52042: data = 8'h05;
      17'd52043: data = 8'h02;
      17'd52044: data = 8'hfe;
      17'd52045: data = 8'hf9;
      17'd52046: data = 8'hf2;
      17'd52047: data = 8'hf1;
      17'd52048: data = 8'hed;
      17'd52049: data = 8'heb;
      17'd52050: data = 8'hf2;
      17'd52051: data = 8'hf6;
      17'd52052: data = 8'hf6;
      17'd52053: data = 8'hf6;
      17'd52054: data = 8'hf4;
      17'd52055: data = 8'hf1;
      17'd52056: data = 8'hf1;
      17'd52057: data = 8'hf1;
      17'd52058: data = 8'hf4;
      17'd52059: data = 8'hfc;
      17'd52060: data = 8'h01;
      17'd52061: data = 8'h06;
      17'd52062: data = 8'h06;
      17'd52063: data = 8'h09;
      17'd52064: data = 8'h0e;
      17'd52065: data = 8'h12;
      17'd52066: data = 8'h13;
      17'd52067: data = 8'h15;
      17'd52068: data = 8'h16;
      17'd52069: data = 8'h16;
      17'd52070: data = 8'h16;
      17'd52071: data = 8'h15;
      17'd52072: data = 8'h0e;
      17'd52073: data = 8'h0a;
      17'd52074: data = 8'h06;
      17'd52075: data = 8'h02;
      17'd52076: data = 8'h00;
      17'd52077: data = 8'hfd;
      17'd52078: data = 8'hfe;
      17'd52079: data = 8'hfa;
      17'd52080: data = 8'hf2;
      17'd52081: data = 8'hef;
      17'd52082: data = 8'hef;
      17'd52083: data = 8'heb;
      17'd52084: data = 8'he9;
      17'd52085: data = 8'he9;
      17'd52086: data = 8'he4;
      17'd52087: data = 8'he3;
      17'd52088: data = 8'he4;
      17'd52089: data = 8'he7;
      17'd52090: data = 8'hec;
      17'd52091: data = 8'hef;
      17'd52092: data = 8'hf4;
      17'd52093: data = 8'hf9;
      17'd52094: data = 8'hfe;
      17'd52095: data = 8'h04;
      17'd52096: data = 8'h09;
      17'd52097: data = 8'h09;
      17'd52098: data = 8'h06;
      17'd52099: data = 8'h06;
      17'd52100: data = 8'h05;
      17'd52101: data = 8'h05;
      17'd52102: data = 8'h00;
      17'd52103: data = 8'hfa;
      17'd52104: data = 8'hf9;
      17'd52105: data = 8'hf9;
      17'd52106: data = 8'hfa;
      17'd52107: data = 8'hfa;
      17'd52108: data = 8'hfa;
      17'd52109: data = 8'hf6;
      17'd52110: data = 8'hf5;
      17'd52111: data = 8'hf4;
      17'd52112: data = 8'hf5;
      17'd52113: data = 8'hf9;
      17'd52114: data = 8'hf6;
      17'd52115: data = 8'hf2;
      17'd52116: data = 8'hef;
      17'd52117: data = 8'hef;
      17'd52118: data = 8'hef;
      17'd52119: data = 8'hf1;
      17'd52120: data = 8'hf4;
      17'd52121: data = 8'hef;
      17'd52122: data = 8'heb;
      17'd52123: data = 8'hef;
      17'd52124: data = 8'hf1;
      17'd52125: data = 8'hf2;
      17'd52126: data = 8'hf4;
      17'd52127: data = 8'hf2;
      17'd52128: data = 8'hef;
      17'd52129: data = 8'hf2;
      17'd52130: data = 8'hf2;
      17'd52131: data = 8'hf6;
      17'd52132: data = 8'hf6;
      17'd52133: data = 8'hfc;
      17'd52134: data = 8'hfc;
      17'd52135: data = 8'hfc;
      17'd52136: data = 8'h01;
      17'd52137: data = 8'h04;
      17'd52138: data = 8'h02;
      17'd52139: data = 8'h02;
      17'd52140: data = 8'h02;
      17'd52141: data = 8'h02;
      17'd52142: data = 8'h04;
      17'd52143: data = 8'h02;
      17'd52144: data = 8'h00;
      17'd52145: data = 8'hfe;
      17'd52146: data = 8'hfd;
      17'd52147: data = 8'hfe;
      17'd52148: data = 8'h01;
      17'd52149: data = 8'h02;
      17'd52150: data = 8'h02;
      17'd52151: data = 8'h05;
      17'd52152: data = 8'h0a;
      17'd52153: data = 8'h0c;
      17'd52154: data = 8'h0c;
      17'd52155: data = 8'h0a;
      17'd52156: data = 8'h05;
      17'd52157: data = 8'h09;
      17'd52158: data = 8'h09;
      17'd52159: data = 8'h0a;
      17'd52160: data = 8'h0c;
      17'd52161: data = 8'h09;
      17'd52162: data = 8'h06;
      17'd52163: data = 8'h04;
      17'd52164: data = 8'h02;
      17'd52165: data = 8'h02;
      17'd52166: data = 8'hfe;
      17'd52167: data = 8'h02;
      17'd52168: data = 8'h02;
      17'd52169: data = 8'h00;
      17'd52170: data = 8'h01;
      17'd52171: data = 8'hfd;
      17'd52172: data = 8'hf9;
      17'd52173: data = 8'hfa;
      17'd52174: data = 8'hfa;
      17'd52175: data = 8'hfa;
      17'd52176: data = 8'hfc;
      17'd52177: data = 8'hfa;
      17'd52178: data = 8'hf6;
      17'd52179: data = 8'hfc;
      17'd52180: data = 8'h01;
      17'd52181: data = 8'h02;
      17'd52182: data = 8'h06;
      17'd52183: data = 8'h0a;
      17'd52184: data = 8'h0c;
      17'd52185: data = 8'h11;
      17'd52186: data = 8'h12;
      17'd52187: data = 8'h0a;
      17'd52188: data = 8'h0c;
      17'd52189: data = 8'h11;
      17'd52190: data = 8'h19;
      17'd52191: data = 8'h1c;
      17'd52192: data = 8'h1b;
      17'd52193: data = 8'h22;
      17'd52194: data = 8'h19;
      17'd52195: data = 8'h19;
      17'd52196: data = 8'h1e;
      17'd52197: data = 8'h0e;
      17'd52198: data = 8'h11;
      17'd52199: data = 8'h0a;
      17'd52200: data = 8'hfa;
      17'd52201: data = 8'hfa;
      17'd52202: data = 8'hf9;
      17'd52203: data = 8'hf6;
      17'd52204: data = 8'hfa;
      17'd52205: data = 8'h04;
      17'd52206: data = 8'h0e;
      17'd52207: data = 8'h05;
      17'd52208: data = 8'hf1;
      17'd52209: data = 8'hdc;
      17'd52210: data = 8'hbd;
      17'd52211: data = 8'hc2;
      17'd52212: data = 8'he0;
      17'd52213: data = 8'hf9;
      17'd52214: data = 8'h1a;
      17'd52215: data = 8'h1f;
      17'd52216: data = 8'h2b;
      17'd52217: data = 8'h24;
      17'd52218: data = 8'h22;
      17'd52219: data = 8'h2f;
      17'd52220: data = 8'h2d;
      17'd52221: data = 8'h35;
      17'd52222: data = 8'h39;
      17'd52223: data = 8'h3a;
      17'd52224: data = 8'h39;
      17'd52225: data = 8'h34;
      17'd52226: data = 8'h1c;
      17'd52227: data = 8'hf5;
      17'd52228: data = 8'hc0;
      17'd52229: data = 8'ha1;
      17'd52230: data = 8'h94;
      17'd52231: data = 8'hae;
      17'd52232: data = 8'hdc;
      17'd52233: data = 8'h06;
      17'd52234: data = 8'h1b;
      17'd52235: data = 8'h0d;
      17'd52236: data = 8'hef;
      17'd52237: data = 8'hd8;
      17'd52238: data = 8'he4;
      17'd52239: data = 8'h04;
      17'd52240: data = 8'h3d;
      17'd52241: data = 8'h64;
      17'd52242: data = 8'h65;
      17'd52243: data = 8'h53;
      17'd52244: data = 8'h27;
      17'd52245: data = 8'hfc;
      17'd52246: data = 8'he4;
      17'd52247: data = 8'he4;
      17'd52248: data = 8'hec;
      17'd52249: data = 8'hf4;
      17'd52250: data = 8'hf2;
      17'd52251: data = 8'hdc;
      17'd52252: data = 8'hbd;
      17'd52253: data = 8'hb3;
      17'd52254: data = 8'hb3;
      17'd52255: data = 8'hbd;
      17'd52256: data = 8'hca;
      17'd52257: data = 8'hdb;
      17'd52258: data = 8'heb;
      17'd52259: data = 8'h00;
      17'd52260: data = 8'h22;
      17'd52261: data = 8'h36;
      17'd52262: data = 8'h42;
      17'd52263: data = 8'h34;
      17'd52264: data = 8'h1f;
      17'd52265: data = 8'h05;
      17'd52266: data = 8'hfe;
      17'd52267: data = 8'h0a;
      17'd52268: data = 8'h16;
      17'd52269: data = 8'h19;
      17'd52270: data = 8'h01;
      17'd52271: data = 8'he3;
      17'd52272: data = 8'hbd;
      17'd52273: data = 8'ha2;
      17'd52274: data = 8'h9a;
      17'd52275: data = 8'ha8;
      17'd52276: data = 8'hbd;
      17'd52277: data = 8'hdb;
      17'd52278: data = 8'hf2;
      17'd52279: data = 8'hf9;
      17'd52280: data = 8'hed;
      17'd52281: data = 8'he9;
      17'd52282: data = 8'hed;
      17'd52283: data = 8'hfd;
      17'd52284: data = 8'h16;
      17'd52285: data = 8'h31;
      17'd52286: data = 8'h3c;
      17'd52287: data = 8'h34;
      17'd52288: data = 8'h2c;
      17'd52289: data = 8'h1f;
      17'd52290: data = 8'h13;
      17'd52291: data = 8'h0c;
      17'd52292: data = 8'h09;
      17'd52293: data = 8'h06;
      17'd52294: data = 8'h02;
      17'd52295: data = 8'h04;
      17'd52296: data = 8'h09;
      17'd52297: data = 8'h06;
      17'd52298: data = 8'h04;
      17'd52299: data = 8'h06;
      17'd52300: data = 8'h05;
      17'd52301: data = 8'h06;
      17'd52302: data = 8'h0e;
      17'd52303: data = 8'h1a;
      17'd52304: data = 8'h22;
      17'd52305: data = 8'h29;
      17'd52306: data = 8'h2c;
      17'd52307: data = 8'h29;
      17'd52308: data = 8'h1f;
      17'd52309: data = 8'h12;
      17'd52310: data = 8'h06;
      17'd52311: data = 8'hfc;
      17'd52312: data = 8'hf2;
      17'd52313: data = 8'hec;
      17'd52314: data = 8'he5;
      17'd52315: data = 8'hdb;
      17'd52316: data = 8'hd1;
      17'd52317: data = 8'hcb;
      17'd52318: data = 8'hc5;
      17'd52319: data = 8'hc5;
      17'd52320: data = 8'hcb;
      17'd52321: data = 8'hd5;
      17'd52322: data = 8'hd8;
      17'd52323: data = 8'he0;
      17'd52324: data = 8'hec;
      17'd52325: data = 8'hf1;
      17'd52326: data = 8'hf9;
      17'd52327: data = 8'hfe;
      17'd52328: data = 8'h06;
      17'd52329: data = 8'h0c;
      17'd52330: data = 8'h09;
      17'd52331: data = 8'h0a;
      17'd52332: data = 8'h0a;
      17'd52333: data = 8'h0a;
      17'd52334: data = 8'h0a;
      17'd52335: data = 8'h0e;
      17'd52336: data = 8'h11;
      17'd52337: data = 8'h0a;
      17'd52338: data = 8'h05;
      17'd52339: data = 8'h06;
      17'd52340: data = 8'h04;
      17'd52341: data = 8'h02;
      17'd52342: data = 8'h09;
      17'd52343: data = 8'h09;
      17'd52344: data = 8'h05;
      17'd52345: data = 8'h05;
      17'd52346: data = 8'h05;
      17'd52347: data = 8'h02;
      17'd52348: data = 8'hfe;
      17'd52349: data = 8'hfe;
      17'd52350: data = 8'hfc;
      17'd52351: data = 8'hf6;
      17'd52352: data = 8'hf9;
      17'd52353: data = 8'hfa;
      17'd52354: data = 8'hf6;
      17'd52355: data = 8'hf1;
      17'd52356: data = 8'heb;
      17'd52357: data = 8'he5;
      17'd52358: data = 8'he2;
      17'd52359: data = 8'hde;
      17'd52360: data = 8'he2;
      17'd52361: data = 8'he4;
      17'd52362: data = 8'he5;
      17'd52363: data = 8'he9;
      17'd52364: data = 8'hec;
      17'd52365: data = 8'heb;
      17'd52366: data = 8'heb;
      17'd52367: data = 8'hec;
      17'd52368: data = 8'hec;
      17'd52369: data = 8'hed;
      17'd52370: data = 8'hf6;
      17'd52371: data = 8'hfd;
      17'd52372: data = 8'hfa;
      17'd52373: data = 8'hf1;
      17'd52374: data = 8'hed;
      17'd52375: data = 8'hed;
      17'd52376: data = 8'hef;
      17'd52377: data = 8'hf6;
      17'd52378: data = 8'hfe;
      17'd52379: data = 8'h04;
      17'd52380: data = 8'h09;
      17'd52381: data = 8'h06;
      17'd52382: data = 8'h06;
      17'd52383: data = 8'h06;
      17'd52384: data = 8'h06;
      17'd52385: data = 8'h0d;
      17'd52386: data = 8'h11;
      17'd52387: data = 8'h11;
      17'd52388: data = 8'h12;
      17'd52389: data = 8'h11;
      17'd52390: data = 8'h0c;
      17'd52391: data = 8'h04;
      17'd52392: data = 8'hfa;
      17'd52393: data = 8'hf1;
      17'd52394: data = 8'hed;
      17'd52395: data = 8'hf1;
      17'd52396: data = 8'hf9;
      17'd52397: data = 8'h04;
      17'd52398: data = 8'h09;
      17'd52399: data = 8'h06;
      17'd52400: data = 8'hfe;
      17'd52401: data = 8'hfc;
      17'd52402: data = 8'hfe;
      17'd52403: data = 8'h02;
      17'd52404: data = 8'h11;
      17'd52405: data = 8'h1b;
      17'd52406: data = 8'h1b;
      17'd52407: data = 8'h19;
      17'd52408: data = 8'h0e;
      17'd52409: data = 8'h05;
      17'd52410: data = 8'h01;
      17'd52411: data = 8'h01;
      17'd52412: data = 8'h05;
      17'd52413: data = 8'h09;
      17'd52414: data = 8'h09;
      17'd52415: data = 8'h06;
      17'd52416: data = 8'h01;
      17'd52417: data = 8'hf9;
      17'd52418: data = 8'hf9;
      17'd52419: data = 8'hf6;
      17'd52420: data = 8'hfa;
      17'd52421: data = 8'h00;
      17'd52422: data = 8'h00;
      17'd52423: data = 8'h05;
      17'd52424: data = 8'h05;
      17'd52425: data = 8'h04;
      17'd52426: data = 8'h0a;
      17'd52427: data = 8'h0c;
      17'd52428: data = 8'h0a;
      17'd52429: data = 8'h11;
      17'd52430: data = 8'h0d;
      17'd52431: data = 8'h12;
      17'd52432: data = 8'h13;
      17'd52433: data = 8'h0e;
      17'd52434: data = 8'h0e;
      17'd52435: data = 8'h02;
      17'd52436: data = 8'h02;
      17'd52437: data = 8'hfc;
      17'd52438: data = 8'hf2;
      17'd52439: data = 8'hfa;
      17'd52440: data = 8'hf6;
      17'd52441: data = 8'hfa;
      17'd52442: data = 8'hfd;
      17'd52443: data = 8'hfa;
      17'd52444: data = 8'h01;
      17'd52445: data = 8'hfa;
      17'd52446: data = 8'hf9;
      17'd52447: data = 8'h02;
      17'd52448: data = 8'h09;
      17'd52449: data = 8'h12;
      17'd52450: data = 8'h15;
      17'd52451: data = 8'h13;
      17'd52452: data = 8'h12;
      17'd52453: data = 8'h0c;
      17'd52454: data = 8'h0a;
      17'd52455: data = 8'h0d;
      17'd52456: data = 8'h0c;
      17'd52457: data = 8'h09;
      17'd52458: data = 8'h06;
      17'd52459: data = 8'h06;
      17'd52460: data = 8'h05;
      17'd52461: data = 8'hfd;
      17'd52462: data = 8'hf6;
      17'd52463: data = 8'hf4;
      17'd52464: data = 8'hf2;
      17'd52465: data = 8'hf9;
      17'd52466: data = 8'h00;
      17'd52467: data = 8'h04;
      17'd52468: data = 8'h04;
      17'd52469: data = 8'h01;
      17'd52470: data = 8'h00;
      17'd52471: data = 8'h04;
      17'd52472: data = 8'h06;
      17'd52473: data = 8'h09;
      17'd52474: data = 8'h0d;
      17'd52475: data = 8'h13;
      17'd52476: data = 8'h16;
      17'd52477: data = 8'h1a;
      17'd52478: data = 8'h1f;
      17'd52479: data = 8'h1e;
      17'd52480: data = 8'h19;
      17'd52481: data = 8'h12;
      17'd52482: data = 8'h12;
      17'd52483: data = 8'h13;
      17'd52484: data = 8'h19;
      17'd52485: data = 8'h19;
      17'd52486: data = 8'h15;
      17'd52487: data = 8'h13;
      17'd52488: data = 8'h0a;
      17'd52489: data = 8'h04;
      17'd52490: data = 8'h00;
      17'd52491: data = 8'hfe;
      17'd52492: data = 8'hfe;
      17'd52493: data = 8'h01;
      17'd52494: data = 8'h06;
      17'd52495: data = 8'h01;
      17'd52496: data = 8'hf4;
      17'd52497: data = 8'hed;
      17'd52498: data = 8'he4;
      17'd52499: data = 8'he5;
      17'd52500: data = 8'he3;
      17'd52501: data = 8'he5;
      17'd52502: data = 8'he5;
      17'd52503: data = 8'hdc;
      17'd52504: data = 8'hdb;
      17'd52505: data = 8'hda;
      17'd52506: data = 8'hdb;
      17'd52507: data = 8'hdb;
      17'd52508: data = 8'hd6;
      17'd52509: data = 8'hd6;
      17'd52510: data = 8'hd8;
      17'd52511: data = 8'hd6;
      17'd52512: data = 8'hdc;
      17'd52513: data = 8'he2;
      17'd52514: data = 8'he7;
      17'd52515: data = 8'hed;
      17'd52516: data = 8'hf4;
      17'd52517: data = 8'hfe;
      17'd52518: data = 8'hfc;
      17'd52519: data = 8'hf5;
      17'd52520: data = 8'hf4;
      17'd52521: data = 8'hf9;
      17'd52522: data = 8'h02;
      17'd52523: data = 8'h0c;
      17'd52524: data = 8'h11;
      17'd52525: data = 8'h11;
      17'd52526: data = 8'h0e;
      17'd52527: data = 8'h12;
      17'd52528: data = 8'h15;
      17'd52529: data = 8'h1a;
      17'd52530: data = 8'h1a;
      17'd52531: data = 8'h16;
      17'd52532: data = 8'h16;
      17'd52533: data = 8'h1c;
      17'd52534: data = 8'h24;
      17'd52535: data = 8'h24;
      17'd52536: data = 8'h23;
      17'd52537: data = 8'h1f;
      17'd52538: data = 8'h1a;
      17'd52539: data = 8'h15;
      17'd52540: data = 8'h11;
      17'd52541: data = 8'h13;
      17'd52542: data = 8'h1a;
      17'd52543: data = 8'h19;
      17'd52544: data = 8'h19;
      17'd52545: data = 8'h1a;
      17'd52546: data = 8'h12;
      17'd52547: data = 8'h09;
      17'd52548: data = 8'hfd;
      17'd52549: data = 8'hf9;
      17'd52550: data = 8'hf6;
      17'd52551: data = 8'hfc;
      17'd52552: data = 8'h02;
      17'd52553: data = 8'h01;
      17'd52554: data = 8'hf6;
      17'd52555: data = 8'hef;
      17'd52556: data = 8'he7;
      17'd52557: data = 8'he5;
      17'd52558: data = 8'he9;
      17'd52559: data = 8'he9;
      17'd52560: data = 8'hed;
      17'd52561: data = 8'hf2;
      17'd52562: data = 8'hf1;
      17'd52563: data = 8'heb;
      17'd52564: data = 8'he3;
      17'd52565: data = 8'hda;
      17'd52566: data = 8'hd3;
      17'd52567: data = 8'hd1;
      17'd52568: data = 8'hd5;
      17'd52569: data = 8'he0;
      17'd52570: data = 8'he5;
      17'd52571: data = 8'he4;
      17'd52572: data = 8'he3;
      17'd52573: data = 8'he7;
      17'd52574: data = 8'he4;
      17'd52575: data = 8'he5;
      17'd52576: data = 8'hed;
      17'd52577: data = 8'hf1;
      17'd52578: data = 8'hfa;
      17'd52579: data = 8'h02;
      17'd52580: data = 8'h0a;
      17'd52581: data = 8'h0e;
      17'd52582: data = 8'h0a;
      17'd52583: data = 8'h05;
      17'd52584: data = 8'h02;
      17'd52585: data = 8'h04;
      17'd52586: data = 8'h09;
      17'd52587: data = 8'h0d;
      17'd52588: data = 8'h11;
      17'd52589: data = 8'h12;
      17'd52590: data = 8'h0e;
      17'd52591: data = 8'h0c;
      17'd52592: data = 8'h05;
      17'd52593: data = 8'h01;
      17'd52594: data = 8'hfd;
      17'd52595: data = 8'hfd;
      17'd52596: data = 8'h02;
      17'd52597: data = 8'h09;
      17'd52598: data = 8'h0a;
      17'd52599: data = 8'h04;
      17'd52600: data = 8'hfd;
      17'd52601: data = 8'hf6;
      17'd52602: data = 8'hf1;
      17'd52603: data = 8'hed;
      17'd52604: data = 8'hf1;
      17'd52605: data = 8'hf2;
      17'd52606: data = 8'hf1;
      17'd52607: data = 8'hef;
      17'd52608: data = 8'heb;
      17'd52609: data = 8'he4;
      17'd52610: data = 8'hdc;
      17'd52611: data = 8'hd6;
      17'd52612: data = 8'hd8;
      17'd52613: data = 8'hdc;
      17'd52614: data = 8'he3;
      17'd52615: data = 8'he7;
      17'd52616: data = 8'heb;
      17'd52617: data = 8'he7;
      17'd52618: data = 8'he3;
      17'd52619: data = 8'he2;
      17'd52620: data = 8'he4;
      17'd52621: data = 8'heb;
      17'd52622: data = 8'hed;
      17'd52623: data = 8'hf2;
      17'd52624: data = 8'hf6;
      17'd52625: data = 8'hf6;
      17'd52626: data = 8'hf5;
      17'd52627: data = 8'hf1;
      17'd52628: data = 8'hef;
      17'd52629: data = 8'hf1;
      17'd52630: data = 8'hf4;
      17'd52631: data = 8'hfa;
      17'd52632: data = 8'h01;
      17'd52633: data = 8'h04;
      17'd52634: data = 8'h00;
      17'd52635: data = 8'hfe;
      17'd52636: data = 8'h02;
      17'd52637: data = 8'h04;
      17'd52638: data = 8'h0c;
      17'd52639: data = 8'h12;
      17'd52640: data = 8'h15;
      17'd52641: data = 8'h16;
      17'd52642: data = 8'h15;
      17'd52643: data = 8'h1a;
      17'd52644: data = 8'h16;
      17'd52645: data = 8'h13;
      17'd52646: data = 8'h13;
      17'd52647: data = 8'h15;
      17'd52648: data = 8'h1a;
      17'd52649: data = 8'h1c;
      17'd52650: data = 8'h1e;
      17'd52651: data = 8'h1a;
      17'd52652: data = 8'h13;
      17'd52653: data = 8'h12;
      17'd52654: data = 8'h13;
      17'd52655: data = 8'h13;
      17'd52656: data = 8'h0e;
      17'd52657: data = 8'h0d;
      17'd52658: data = 8'h0c;
      17'd52659: data = 8'h09;
      17'd52660: data = 8'h02;
      17'd52661: data = 8'hfc;
      17'd52662: data = 8'hf4;
      17'd52663: data = 8'hed;
      17'd52664: data = 8'heb;
      17'd52665: data = 8'hf1;
      17'd52666: data = 8'hf2;
      17'd52667: data = 8'hf1;
      17'd52668: data = 8'hf1;
      17'd52669: data = 8'hf1;
      17'd52670: data = 8'hfa;
      17'd52671: data = 8'hfc;
      17'd52672: data = 8'h02;
      17'd52673: data = 8'h06;
      17'd52674: data = 8'h05;
      17'd52675: data = 8'h09;
      17'd52676: data = 8'h09;
      17'd52677: data = 8'h0c;
      17'd52678: data = 8'h05;
      17'd52679: data = 8'hfd;
      17'd52680: data = 8'h00;
      17'd52681: data = 8'h05;
      17'd52682: data = 8'h09;
      17'd52683: data = 8'h0d;
      17'd52684: data = 8'h0a;
      17'd52685: data = 8'h09;
      17'd52686: data = 8'h09;
      17'd52687: data = 8'h06;
      17'd52688: data = 8'h0e;
      17'd52689: data = 8'h15;
      17'd52690: data = 8'h13;
      17'd52691: data = 8'h1a;
      17'd52692: data = 8'h1a;
      17'd52693: data = 8'h19;
      17'd52694: data = 8'h16;
      17'd52695: data = 8'h0c;
      17'd52696: data = 8'h0a;
      17'd52697: data = 8'h0e;
      17'd52698: data = 8'h12;
      17'd52699: data = 8'h16;
      17'd52700: data = 8'h1c;
      17'd52701: data = 8'h19;
      17'd52702: data = 8'h16;
      17'd52703: data = 8'h11;
      17'd52704: data = 8'h0a;
      17'd52705: data = 8'h0c;
      17'd52706: data = 8'h05;
      17'd52707: data = 8'h00;
      17'd52708: data = 8'hfc;
      17'd52709: data = 8'hfa;
      17'd52710: data = 8'hf4;
      17'd52711: data = 8'hed;
      17'd52712: data = 8'hef;
      17'd52713: data = 8'hf1;
      17'd52714: data = 8'hf1;
      17'd52715: data = 8'hf1;
      17'd52716: data = 8'hf6;
      17'd52717: data = 8'h01;
      17'd52718: data = 8'h04;
      17'd52719: data = 8'h09;
      17'd52720: data = 8'h11;
      17'd52721: data = 8'h1a;
      17'd52722: data = 8'h1f;
      17'd52723: data = 8'h1e;
      17'd52724: data = 8'h1e;
      17'd52725: data = 8'h1f;
      17'd52726: data = 8'h1e;
      17'd52727: data = 8'h1b;
      17'd52728: data = 8'h1c;
      17'd52729: data = 8'h1b;
      17'd52730: data = 8'h13;
      17'd52731: data = 8'h09;
      17'd52732: data = 8'h0a;
      17'd52733: data = 8'h0c;
      17'd52734: data = 8'h05;
      17'd52735: data = 8'h02;
      17'd52736: data = 8'h06;
      17'd52737: data = 8'h0a;
      17'd52738: data = 8'h06;
      17'd52739: data = 8'h0a;
      17'd52740: data = 8'h0d;
      17'd52741: data = 8'h0e;
      17'd52742: data = 8'h05;
      17'd52743: data = 8'h02;
      17'd52744: data = 8'h09;
      17'd52745: data = 8'h06;
      17'd52746: data = 8'h04;
      17'd52747: data = 8'h00;
      17'd52748: data = 8'hfe;
      17'd52749: data = 8'hfa;
      17'd52750: data = 8'hf1;
      17'd52751: data = 8'heb;
      17'd52752: data = 8'he9;
      17'd52753: data = 8'he4;
      17'd52754: data = 8'he2;
      17'd52755: data = 8'hde;
      17'd52756: data = 8'hdc;
      17'd52757: data = 8'hdc;
      17'd52758: data = 8'hd8;
      17'd52759: data = 8'hd1;
      17'd52760: data = 8'hd1;
      17'd52761: data = 8'hd3;
      17'd52762: data = 8'hd5;
      17'd52763: data = 8'hda;
      17'd52764: data = 8'he3;
      17'd52765: data = 8'he9;
      17'd52766: data = 8'he3;
      17'd52767: data = 8'he3;
      17'd52768: data = 8'he9;
      17'd52769: data = 8'hed;
      17'd52770: data = 8'hed;
      17'd52771: data = 8'hed;
      17'd52772: data = 8'hf4;
      17'd52773: data = 8'hf9;
      17'd52774: data = 8'hf6;
      17'd52775: data = 8'hf6;
      17'd52776: data = 8'hfd;
      17'd52777: data = 8'hfe;
      17'd52778: data = 8'hfd;
      17'd52779: data = 8'hfd;
      17'd52780: data = 8'h02;
      17'd52781: data = 8'h0a;
      17'd52782: data = 8'h0d;
      17'd52783: data = 8'h11;
      17'd52784: data = 8'h13;
      17'd52785: data = 8'h16;
      17'd52786: data = 8'h15;
      17'd52787: data = 8'h12;
      17'd52788: data = 8'h1a;
      17'd52789: data = 8'h1f;
      17'd52790: data = 8'h1f;
      17'd52791: data = 8'h22;
      17'd52792: data = 8'h26;
      17'd52793: data = 8'h24;
      17'd52794: data = 8'h1f;
      17'd52795: data = 8'h1c;
      17'd52796: data = 8'h1e;
      17'd52797: data = 8'h1c;
      17'd52798: data = 8'h1c;
      17'd52799: data = 8'h1b;
      17'd52800: data = 8'h19;
      17'd52801: data = 8'h16;
      17'd52802: data = 8'h12;
      17'd52803: data = 8'h0c;
      17'd52804: data = 8'h06;
      17'd52805: data = 8'h04;
      17'd52806: data = 8'hfe;
      17'd52807: data = 8'hfc;
      17'd52808: data = 8'hfa;
      17'd52809: data = 8'hf6;
      17'd52810: data = 8'hf2;
      17'd52811: data = 8'hec;
      17'd52812: data = 8'he9;
      17'd52813: data = 8'he9;
      17'd52814: data = 8'he7;
      17'd52815: data = 8'he5;
      17'd52816: data = 8'he7;
      17'd52817: data = 8'he7;
      17'd52818: data = 8'he5;
      17'd52819: data = 8'he3;
      17'd52820: data = 8'he0;
      17'd52821: data = 8'he0;
      17'd52822: data = 8'hde;
      17'd52823: data = 8'hdc;
      17'd52824: data = 8'hde;
      17'd52825: data = 8'he0;
      17'd52826: data = 8'he2;
      17'd52827: data = 8'he0;
      17'd52828: data = 8'hdc;
      17'd52829: data = 8'hdc;
      17'd52830: data = 8'hdc;
      17'd52831: data = 8'he0;
      17'd52832: data = 8'he0;
      17'd52833: data = 8'he2;
      17'd52834: data = 8'he7;
      17'd52835: data = 8'he9;
      17'd52836: data = 8'heb;
      17'd52837: data = 8'hed;
      17'd52838: data = 8'hec;
      17'd52839: data = 8'hec;
      17'd52840: data = 8'hed;
      17'd52841: data = 8'hf2;
      17'd52842: data = 8'hf9;
      17'd52843: data = 8'hf9;
      17'd52844: data = 8'hfe;
      17'd52845: data = 8'h02;
      17'd52846: data = 8'h01;
      17'd52847: data = 8'h00;
      17'd52848: data = 8'h00;
      17'd52849: data = 8'hfe;
      17'd52850: data = 8'hfe;
      17'd52851: data = 8'hfd;
      17'd52852: data = 8'hfe;
      17'd52853: data = 8'h02;
      17'd52854: data = 8'h01;
      17'd52855: data = 8'hfe;
      17'd52856: data = 8'hfe;
      17'd52857: data = 8'hfc;
      17'd52858: data = 8'hfc;
      17'd52859: data = 8'hfd;
      17'd52860: data = 8'hfe;
      17'd52861: data = 8'hfe;
      17'd52862: data = 8'h00;
      17'd52863: data = 8'hfe;
      17'd52864: data = 8'hfd;
      17'd52865: data = 8'hfe;
      17'd52866: data = 8'hfc;
      17'd52867: data = 8'hf9;
      17'd52868: data = 8'hf9;
      17'd52869: data = 8'hfa;
      17'd52870: data = 8'hf9;
      17'd52871: data = 8'hf9;
      17'd52872: data = 8'hf9;
      17'd52873: data = 8'hf6;
      17'd52874: data = 8'hf2;
      17'd52875: data = 8'hf1;
      17'd52876: data = 8'hf1;
      17'd52877: data = 8'hf1;
      17'd52878: data = 8'hf2;
      17'd52879: data = 8'hf4;
      17'd52880: data = 8'hf5;
      17'd52881: data = 8'hf5;
      17'd52882: data = 8'hf5;
      17'd52883: data = 8'hf5;
      17'd52884: data = 8'hf6;
      17'd52885: data = 8'hf6;
      17'd52886: data = 8'hfa;
      17'd52887: data = 8'hfd;
      17'd52888: data = 8'hfd;
      17'd52889: data = 8'hfd;
      17'd52890: data = 8'hfe;
      17'd52891: data = 8'hfe;
      17'd52892: data = 8'h00;
      17'd52893: data = 8'h02;
      17'd52894: data = 8'h04;
      17'd52895: data = 8'h04;
      17'd52896: data = 8'h06;
      17'd52897: data = 8'h0c;
      17'd52898: data = 8'h0a;
      17'd52899: data = 8'h0c;
      17'd52900: data = 8'h0c;
      17'd52901: data = 8'h0c;
      17'd52902: data = 8'h0d;
      17'd52903: data = 8'h11;
      17'd52904: data = 8'h15;
      17'd52905: data = 8'h1a;
      17'd52906: data = 8'h19;
      17'd52907: data = 8'h0c;
      17'd52908: data = 8'h05;
      17'd52909: data = 8'h0a;
      17'd52910: data = 8'h13;
      17'd52911: data = 8'h19;
      17'd52912: data = 8'h1a;
      17'd52913: data = 8'h1b;
      17'd52914: data = 8'h19;
      17'd52915: data = 8'h12;
      17'd52916: data = 8'h13;
      17'd52917: data = 8'h12;
      17'd52918: data = 8'h09;
      17'd52919: data = 8'h09;
      17'd52920: data = 8'h13;
      17'd52921: data = 8'h12;
      17'd52922: data = 8'h09;
      17'd52923: data = 8'h0a;
      17'd52924: data = 8'h09;
      17'd52925: data = 8'h01;
      17'd52926: data = 8'h01;
      17'd52927: data = 8'h09;
      17'd52928: data = 8'h04;
      17'd52929: data = 8'hfd;
      17'd52930: data = 8'h02;
      17'd52931: data = 8'h02;
      17'd52932: data = 8'h04;
      17'd52933: data = 8'h02;
      17'd52934: data = 8'hfd;
      17'd52935: data = 8'hf5;
      17'd52936: data = 8'hf9;
      17'd52937: data = 8'hfe;
      17'd52938: data = 8'hfe;
      17'd52939: data = 8'h01;
      17'd52940: data = 8'h09;
      17'd52941: data = 8'h0c;
      17'd52942: data = 8'h0e;
      17'd52943: data = 8'h0e;
      17'd52944: data = 8'h0c;
      17'd52945: data = 8'h02;
      17'd52946: data = 8'h00;
      17'd52947: data = 8'h09;
      17'd52948: data = 8'h05;
      17'd52949: data = 8'h02;
      17'd52950: data = 8'h02;
      17'd52951: data = 8'h01;
      17'd52952: data = 8'hfe;
      17'd52953: data = 8'hfd;
      17'd52954: data = 8'hfe;
      17'd52955: data = 8'h01;
      17'd52956: data = 8'h05;
      17'd52957: data = 8'h0c;
      17'd52958: data = 8'h15;
      17'd52959: data = 8'h19;
      17'd52960: data = 8'h1f;
      17'd52961: data = 8'h27;
      17'd52962: data = 8'h26;
      17'd52963: data = 8'h29;
      17'd52964: data = 8'h2d;
      17'd52965: data = 8'h29;
      17'd52966: data = 8'h2b;
      17'd52967: data = 8'h2f;
      17'd52968: data = 8'h2c;
      17'd52969: data = 8'h2b;
      17'd52970: data = 8'h26;
      17'd52971: data = 8'h23;
      17'd52972: data = 8'h1a;
      17'd52973: data = 8'h11;
      17'd52974: data = 8'h0a;
      17'd52975: data = 8'h05;
      17'd52976: data = 8'h09;
      17'd52977: data = 8'h0c;
      17'd52978: data = 8'h06;
      17'd52979: data = 8'h06;
      17'd52980: data = 8'h09;
      17'd52981: data = 8'h05;
      17'd52982: data = 8'h04;
      17'd52983: data = 8'h02;
      17'd52984: data = 8'h01;
      17'd52985: data = 8'hfd;
      17'd52986: data = 8'hfd;
      17'd52987: data = 8'hfd;
      17'd52988: data = 8'hfc;
      17'd52989: data = 8'hf6;
      17'd52990: data = 8'hed;
      17'd52991: data = 8'he7;
      17'd52992: data = 8'he2;
      17'd52993: data = 8'hd8;
      17'd52994: data = 8'hd3;
      17'd52995: data = 8'hd6;
      17'd52996: data = 8'hd1;
      17'd52997: data = 8'hce;
      17'd52998: data = 8'hd3;
      17'd52999: data = 8'hd3;
      17'd53000: data = 8'hd3;
      17'd53001: data = 8'hd3;
      17'd53002: data = 8'hd1;
      17'd53003: data = 8'hd2;
      17'd53004: data = 8'hd6;
      17'd53005: data = 8'hdc;
      17'd53006: data = 8'he2;
      17'd53007: data = 8'he3;
      17'd53008: data = 8'he7;
      17'd53009: data = 8'he9;
      17'd53010: data = 8'he9;
      17'd53011: data = 8'heb;
      17'd53012: data = 8'hec;
      17'd53013: data = 8'hed;
      17'd53014: data = 8'hf2;
      17'd53015: data = 8'hf6;
      17'd53016: data = 8'hfa;
      17'd53017: data = 8'hfe;
      17'd53018: data = 8'hfe;
      17'd53019: data = 8'h01;
      17'd53020: data = 8'h05;
      17'd53021: data = 8'h0a;
      17'd53022: data = 8'h13;
      17'd53023: data = 8'h1a;
      17'd53024: data = 8'h1e;
      17'd53025: data = 8'h1e;
      17'd53026: data = 8'h23;
      17'd53027: data = 8'h26;
      17'd53028: data = 8'h26;
      17'd53029: data = 8'h26;
      17'd53030: data = 8'h27;
      17'd53031: data = 8'h27;
      17'd53032: data = 8'h29;
      17'd53033: data = 8'h29;
      17'd53034: data = 8'h27;
      17'd53035: data = 8'h27;
      17'd53036: data = 8'h24;
      17'd53037: data = 8'h1e;
      17'd53038: data = 8'h1f;
      17'd53039: data = 8'h1e;
      17'd53040: data = 8'h1a;
      17'd53041: data = 8'h19;
      17'd53042: data = 8'h13;
      17'd53043: data = 8'h12;
      17'd53044: data = 8'h11;
      17'd53045: data = 8'h0c;
      17'd53046: data = 8'h06;
      17'd53047: data = 8'h05;
      17'd53048: data = 8'h01;
      17'd53049: data = 8'h00;
      17'd53050: data = 8'h00;
      17'd53051: data = 8'hfd;
      17'd53052: data = 8'hf2;
      17'd53053: data = 8'heb;
      17'd53054: data = 8'he9;
      17'd53055: data = 8'he2;
      17'd53056: data = 8'he0;
      17'd53057: data = 8'he2;
      17'd53058: data = 8'hde;
      17'd53059: data = 8'hdc;
      17'd53060: data = 8'hda;
      17'd53061: data = 8'hd8;
      17'd53062: data = 8'hd5;
      17'd53063: data = 8'hd5;
      17'd53064: data = 8'hd8;
      17'd53065: data = 8'hd8;
      17'd53066: data = 8'hdb;
      17'd53067: data = 8'he4;
      17'd53068: data = 8'he5;
      17'd53069: data = 8'hde;
      17'd53070: data = 8'hdc;
      17'd53071: data = 8'hdb;
      17'd53072: data = 8'hdb;
      17'd53073: data = 8'hde;
      17'd53074: data = 8'he2;
      17'd53075: data = 8'he4;
      17'd53076: data = 8'he0;
      17'd53077: data = 8'he2;
      17'd53078: data = 8'he5;
      17'd53079: data = 8'he4;
      17'd53080: data = 8'he2;
      17'd53081: data = 8'he0;
      17'd53082: data = 8'he4;
      17'd53083: data = 8'hed;
      17'd53084: data = 8'hf2;
      17'd53085: data = 8'hfa;
      17'd53086: data = 8'hfc;
      17'd53087: data = 8'hf9;
      17'd53088: data = 8'hfa;
      17'd53089: data = 8'hfe;
      17'd53090: data = 8'h00;
      17'd53091: data = 8'h01;
      17'd53092: data = 8'h02;
      17'd53093: data = 8'h01;
      17'd53094: data = 8'h02;
      17'd53095: data = 8'h05;
      17'd53096: data = 8'h02;
      17'd53097: data = 8'hfe;
      17'd53098: data = 8'hfa;
      17'd53099: data = 8'hfe;
      17'd53100: data = 8'h00;
      17'd53101: data = 8'h01;
      17'd53102: data = 8'h09;
      17'd53103: data = 8'h09;
      17'd53104: data = 8'h04;
      17'd53105: data = 8'hfe;
      17'd53106: data = 8'h00;
      17'd53107: data = 8'h01;
      17'd53108: data = 8'h01;
      17'd53109: data = 8'h05;
      17'd53110: data = 8'h01;
      17'd53111: data = 8'hfa;
      17'd53112: data = 8'hf9;
      17'd53113: data = 8'hfa;
      17'd53114: data = 8'hf2;
      17'd53115: data = 8'heb;
      17'd53116: data = 8'hef;
      17'd53117: data = 8'hf4;
      17'd53118: data = 8'hf4;
      17'd53119: data = 8'hf9;
      17'd53120: data = 8'hf6;
      17'd53121: data = 8'hf2;
      17'd53122: data = 8'hf1;
      17'd53123: data = 8'hef;
      17'd53124: data = 8'hf2;
      17'd53125: data = 8'hf5;
      17'd53126: data = 8'hf6;
      17'd53127: data = 8'hf9;
      17'd53128: data = 8'hf6;
      17'd53129: data = 8'hf6;
      17'd53130: data = 8'hf9;
      17'd53131: data = 8'hf5;
      17'd53132: data = 8'hf2;
      17'd53133: data = 8'hf4;
      17'd53134: data = 8'hfd;
      17'd53135: data = 8'h05;
      17'd53136: data = 8'h0a;
      17'd53137: data = 8'h05;
      17'd53138: data = 8'hfe;
      17'd53139: data = 8'hfe;
      17'd53140: data = 8'h09;
      17'd53141: data = 8'h0c;
      17'd53142: data = 8'h09;
      17'd53143: data = 8'h0a;
      17'd53144: data = 8'h11;
      17'd53145: data = 8'h0d;
      17'd53146: data = 8'h06;
      17'd53147: data = 8'h05;
      17'd53148: data = 8'h04;
      17'd53149: data = 8'h04;
      17'd53150: data = 8'h0d;
      17'd53151: data = 8'h19;
      17'd53152: data = 8'h1b;
      17'd53153: data = 8'h1b;
      17'd53154: data = 8'h19;
      17'd53155: data = 8'h1c;
      17'd53156: data = 8'h1b;
      17'd53157: data = 8'h15;
      17'd53158: data = 8'h16;
      17'd53159: data = 8'h1b;
      17'd53160: data = 8'h1c;
      17'd53161: data = 8'h1b;
      17'd53162: data = 8'h1c;
      17'd53163: data = 8'h1b;
      17'd53164: data = 8'h16;
      17'd53165: data = 8'h0e;
      17'd53166: data = 8'h0e;
      17'd53167: data = 8'h0c;
      17'd53168: data = 8'h0a;
      17'd53169: data = 8'h0c;
      17'd53170: data = 8'h09;
      17'd53171: data = 8'h0a;
      17'd53172: data = 8'h0d;
      17'd53173: data = 8'h05;
      17'd53174: data = 8'h00;
      17'd53175: data = 8'h02;
      17'd53176: data = 8'h00;
      17'd53177: data = 8'hfd;
      17'd53178: data = 8'h01;
      17'd53179: data = 8'h02;
      17'd53180: data = 8'h02;
      17'd53181: data = 8'h0c;
      17'd53182: data = 8'h0d;
      17'd53183: data = 8'h0d;
      17'd53184: data = 8'h06;
      17'd53185: data = 8'hfa;
      17'd53186: data = 8'hfa;
      17'd53187: data = 8'hf4;
      17'd53188: data = 8'hec;
      17'd53189: data = 8'he7;
      17'd53190: data = 8'he9;
      17'd53191: data = 8'hf4;
      17'd53192: data = 8'hed;
      17'd53193: data = 8'hef;
      17'd53194: data = 8'hfd;
      17'd53195: data = 8'hf4;
      17'd53196: data = 8'hf1;
      17'd53197: data = 8'hfc;
      17'd53198: data = 8'h01;
      17'd53199: data = 8'h0e;
      17'd53200: data = 8'h1f;
      17'd53201: data = 8'h2d;
      17'd53202: data = 8'h31;
      17'd53203: data = 8'h31;
      17'd53204: data = 8'h2f;
      17'd53205: data = 8'h23;
      17'd53206: data = 8'h24;
      17'd53207: data = 8'h2d;
      17'd53208: data = 8'h24;
      17'd53209: data = 8'h2b;
      17'd53210: data = 8'h36;
      17'd53211: data = 8'h33;
      17'd53212: data = 8'h2b;
      17'd53213: data = 8'h22;
      17'd53214: data = 8'h1f;
      17'd53215: data = 8'h1a;
      17'd53216: data = 8'h19;
      17'd53217: data = 8'h24;
      17'd53218: data = 8'h27;
      17'd53219: data = 8'h26;
      17'd53220: data = 8'h2b;
      17'd53221: data = 8'h23;
      17'd53222: data = 8'h1f;
      17'd53223: data = 8'h1a;
      17'd53224: data = 8'h0d;
      17'd53225: data = 8'h0d;
      17'd53226: data = 8'h0a;
      17'd53227: data = 8'h0c;
      17'd53228: data = 8'h05;
      17'd53229: data = 8'hfe;
      17'd53230: data = 8'hfa;
      17'd53231: data = 8'heb;
      17'd53232: data = 8'hdc;
      17'd53233: data = 8'hd3;
      17'd53234: data = 8'hd1;
      17'd53235: data = 8'hcd;
      17'd53236: data = 8'hc9;
      17'd53237: data = 8'hcb;
      17'd53238: data = 8'hca;
      17'd53239: data = 8'hc2;
      17'd53240: data = 8'hc4;
      17'd53241: data = 8'hbd;
      17'd53242: data = 8'hbb;
      17'd53243: data = 8'hc0;
      17'd53244: data = 8'hc4;
      17'd53245: data = 8'hca;
      17'd53246: data = 8'hd1;
      17'd53247: data = 8'hd3;
      17'd53248: data = 8'hce;
      17'd53249: data = 8'hc9;
      17'd53250: data = 8'hca;
      17'd53251: data = 8'hcb;
      17'd53252: data = 8'hce;
      17'd53253: data = 8'hdb;
      17'd53254: data = 8'he3;
      17'd53255: data = 8'he7;
      17'd53256: data = 8'hf1;
      17'd53257: data = 8'hf4;
      17'd53258: data = 8'hf6;
      17'd53259: data = 8'hfa;
      17'd53260: data = 8'h01;
      17'd53261: data = 8'h0c;
      17'd53262: data = 8'h16;
      17'd53263: data = 8'h23;
      17'd53264: data = 8'h26;
      17'd53265: data = 8'h2b;
      17'd53266: data = 8'h2c;
      17'd53267: data = 8'h2c;
      17'd53268: data = 8'h2f;
      17'd53269: data = 8'h31;
      17'd53270: data = 8'h34;
      17'd53271: data = 8'h3c;
      17'd53272: data = 8'h3d;
      17'd53273: data = 8'h40;
      17'd53274: data = 8'h40;
      17'd53275: data = 8'h3c;
      17'd53276: data = 8'h3a;
      17'd53277: data = 8'h34;
      17'd53278: data = 8'h33;
      17'd53279: data = 8'h35;
      17'd53280: data = 8'h35;
      17'd53281: data = 8'h36;
      17'd53282: data = 8'h34;
      17'd53283: data = 8'h2b;
      17'd53284: data = 8'h24;
      17'd53285: data = 8'h1b;
      17'd53286: data = 8'h13;
      17'd53287: data = 8'h0d;
      17'd53288: data = 8'h06;
      17'd53289: data = 8'h02;
      17'd53290: data = 8'h00;
      17'd53291: data = 8'hfd;
      17'd53292: data = 8'hf1;
      17'd53293: data = 8'he7;
      17'd53294: data = 8'hdc;
      17'd53295: data = 8'hd3;
      17'd53296: data = 8'hce;
      17'd53297: data = 8'hcd;
      17'd53298: data = 8'hce;
      17'd53299: data = 8'hd1;
      17'd53300: data = 8'hcd;
      17'd53301: data = 8'hc6;
      17'd53302: data = 8'hc5;
      17'd53303: data = 8'hc4;
      17'd53304: data = 8'hc1;
      17'd53305: data = 8'hc0;
      17'd53306: data = 8'hc4;
      17'd53307: data = 8'hc9;
      17'd53308: data = 8'hc9;
      17'd53309: data = 8'hca;
      17'd53310: data = 8'hc5;
      17'd53311: data = 8'hc4;
      17'd53312: data = 8'hc2;
      17'd53313: data = 8'hc4;
      17'd53314: data = 8'hc9;
      17'd53315: data = 8'hd1;
      17'd53316: data = 8'hd8;
      17'd53317: data = 8'he0;
      17'd53318: data = 8'he3;
      17'd53319: data = 8'he3;
      17'd53320: data = 8'he4;
      17'd53321: data = 8'he9;
      17'd53322: data = 8'hec;
      17'd53323: data = 8'hf1;
      17'd53324: data = 8'hfa;
      17'd53325: data = 8'h00;
      17'd53326: data = 8'h01;
      17'd53327: data = 8'h04;
      17'd53328: data = 8'h04;
      17'd53329: data = 8'h04;
      17'd53330: data = 8'h09;
      17'd53331: data = 8'h0a;
      17'd53332: data = 8'h11;
      17'd53333: data = 8'h13;
      17'd53334: data = 8'h15;
      17'd53335: data = 8'h16;
      17'd53336: data = 8'h13;
      17'd53337: data = 8'h13;
      17'd53338: data = 8'h11;
      17'd53339: data = 8'h0d;
      17'd53340: data = 8'h0a;
      17'd53341: data = 8'h0c;
      17'd53342: data = 8'h0d;
      17'd53343: data = 8'h11;
      17'd53344: data = 8'h0e;
      17'd53345: data = 8'h0a;
      17'd53346: data = 8'h09;
      17'd53347: data = 8'h06;
      17'd53348: data = 8'h04;
      17'd53349: data = 8'h00;
      17'd53350: data = 8'hfe;
      17'd53351: data = 8'hfa;
      17'd53352: data = 8'hf5;
      17'd53353: data = 8'hef;
      17'd53354: data = 8'heb;
      17'd53355: data = 8'he7;
      17'd53356: data = 8'he5;
      17'd53357: data = 8'he5;
      17'd53358: data = 8'he7;
      17'd53359: data = 8'he9;
      17'd53360: data = 8'he7;
      17'd53361: data = 8'he9;
      17'd53362: data = 8'he5;
      17'd53363: data = 8'he5;
      17'd53364: data = 8'he5;
      17'd53365: data = 8'he3;
      17'd53366: data = 8'he7;
      17'd53367: data = 8'he7;
      17'd53368: data = 8'he9;
      17'd53369: data = 8'he7;
      17'd53370: data = 8'he5;
      17'd53371: data = 8'he9;
      17'd53372: data = 8'heb;
      17'd53373: data = 8'hed;
      17'd53374: data = 8'hf2;
      17'd53375: data = 8'hf6;
      17'd53376: data = 8'hfa;
      17'd53377: data = 8'h00;
      17'd53378: data = 8'h01;
      17'd53379: data = 8'h00;
      17'd53380: data = 8'h05;
      17'd53381: data = 8'h05;
      17'd53382: data = 8'h06;
      17'd53383: data = 8'h0d;
      17'd53384: data = 8'h13;
      17'd53385: data = 8'h16;
      17'd53386: data = 8'h15;
      17'd53387: data = 8'h19;
      17'd53388: data = 8'h16;
      17'd53389: data = 8'h16;
      17'd53390: data = 8'h1c;
      17'd53391: data = 8'h22;
      17'd53392: data = 8'h22;
      17'd53393: data = 8'h24;
      17'd53394: data = 8'h2c;
      17'd53395: data = 8'h2b;
      17'd53396: data = 8'h23;
      17'd53397: data = 8'h24;
      17'd53398: data = 8'h1e;
      17'd53399: data = 8'h1b;
      17'd53400: data = 8'h1e;
      17'd53401: data = 8'h1b;
      17'd53402: data = 8'h1b;
      17'd53403: data = 8'h1a;
      17'd53404: data = 8'h16;
      17'd53405: data = 8'h11;
      17'd53406: data = 8'h0d;
      17'd53407: data = 8'h0d;
      17'd53408: data = 8'h0a;
      17'd53409: data = 8'h05;
      17'd53410: data = 8'h09;
      17'd53411: data = 8'h09;
      17'd53412: data = 8'h02;
      17'd53413: data = 8'hfe;
      17'd53414: data = 8'h00;
      17'd53415: data = 8'hfe;
      17'd53416: data = 8'hfe;
      17'd53417: data = 8'hfa;
      17'd53418: data = 8'hfd;
      17'd53419: data = 8'hfe;
      17'd53420: data = 8'hfe;
      17'd53421: data = 8'hfe;
      17'd53422: data = 8'hfc;
      17'd53423: data = 8'hfe;
      17'd53424: data = 8'hfe;
      17'd53425: data = 8'h01;
      17'd53426: data = 8'hfe;
      17'd53427: data = 8'hf6;
      17'd53428: data = 8'hf4;
      17'd53429: data = 8'he9;
      17'd53430: data = 8'he7;
      17'd53431: data = 8'hec;
      17'd53432: data = 8'hef;
      17'd53433: data = 8'hf6;
      17'd53434: data = 8'hfa;
      17'd53435: data = 8'hfa;
      17'd53436: data = 8'hfe;
      17'd53437: data = 8'h00;
      17'd53438: data = 8'h06;
      17'd53439: data = 8'h0d;
      17'd53440: data = 8'h16;
      17'd53441: data = 8'h2c;
      17'd53442: data = 8'h33;
      17'd53443: data = 8'h34;
      17'd53444: data = 8'h35;
      17'd53445: data = 8'h31;
      17'd53446: data = 8'h2b;
      17'd53447: data = 8'h26;
      17'd53448: data = 8'h2c;
      17'd53449: data = 8'h2d;
      17'd53450: data = 8'h2b;
      17'd53451: data = 8'h2c;
      17'd53452: data = 8'h2b;
      17'd53453: data = 8'h23;
      17'd53454: data = 8'h1b;
      17'd53455: data = 8'h19;
      17'd53456: data = 8'h16;
      17'd53457: data = 8'h15;
      17'd53458: data = 8'h1c;
      17'd53459: data = 8'h26;
      17'd53460: data = 8'h29;
      17'd53461: data = 8'h27;
      17'd53462: data = 8'h22;
      17'd53463: data = 8'h1c;
      17'd53464: data = 8'h16;
      17'd53465: data = 8'h0e;
      17'd53466: data = 8'h0d;
      17'd53467: data = 8'h06;
      17'd53468: data = 8'h04;
      17'd53469: data = 8'h01;
      17'd53470: data = 8'hf6;
      17'd53471: data = 8'hef;
      17'd53472: data = 8'he4;
      17'd53473: data = 8'hd6;
      17'd53474: data = 8'hd1;
      17'd53475: data = 8'hcd;
      17'd53476: data = 8'hce;
      17'd53477: data = 8'hd3;
      17'd53478: data = 8'hd3;
      17'd53479: data = 8'hd3;
      17'd53480: data = 8'hce;
      17'd53481: data = 8'hca;
      17'd53482: data = 8'hc5;
      17'd53483: data = 8'hc2;
      17'd53484: data = 8'hc6;
      17'd53485: data = 8'hcd;
      17'd53486: data = 8'hd1;
      17'd53487: data = 8'hd5;
      17'd53488: data = 8'hd5;
      17'd53489: data = 8'hd3;
      17'd53490: data = 8'hce;
      17'd53491: data = 8'hcb;
      17'd53492: data = 8'hd2;
      17'd53493: data = 8'hd3;
      17'd53494: data = 8'hda;
      17'd53495: data = 8'he5;
      17'd53496: data = 8'hed;
      17'd53497: data = 8'hed;
      17'd53498: data = 8'hf4;
      17'd53499: data = 8'hf6;
      17'd53500: data = 8'hfd;
      17'd53501: data = 8'h02;
      17'd53502: data = 8'h0a;
      17'd53503: data = 8'h1a;
      17'd53504: data = 8'h23;
      17'd53505: data = 8'h27;
      17'd53506: data = 8'h2c;
      17'd53507: data = 8'h2c;
      17'd53508: data = 8'h29;
      17'd53509: data = 8'h29;
      17'd53510: data = 8'h2b;
      17'd53511: data = 8'h2d;
      17'd53512: data = 8'h34;
      17'd53513: data = 8'h35;
      17'd53514: data = 8'h35;
      17'd53515: data = 8'h33;
      17'd53516: data = 8'h31;
      17'd53517: data = 8'h33;
      17'd53518: data = 8'h33;
      17'd53519: data = 8'h31;
      17'd53520: data = 8'h34;
      17'd53521: data = 8'h35;
      17'd53522: data = 8'h36;
      17'd53523: data = 8'h33;
      17'd53524: data = 8'h29;
      17'd53525: data = 8'h23;
      17'd53526: data = 8'h19;
      17'd53527: data = 8'h11;
      17'd53528: data = 8'h0e;
      17'd53529: data = 8'h0c;
      17'd53530: data = 8'h06;
      17'd53531: data = 8'h04;
      17'd53532: data = 8'hfc;
      17'd53533: data = 8'hf5;
      17'd53534: data = 8'hec;
      17'd53535: data = 8'he3;
      17'd53536: data = 8'hdb;
      17'd53537: data = 8'hda;
      17'd53538: data = 8'hdc;
      17'd53539: data = 8'hda;
      17'd53540: data = 8'hda;
      17'd53541: data = 8'hda;
      17'd53542: data = 8'hd2;
      17'd53543: data = 8'hcb;
      17'd53544: data = 8'hc6;
      17'd53545: data = 8'hc2;
      17'd53546: data = 8'hc4;
      17'd53547: data = 8'hc9;
      17'd53548: data = 8'hcb;
      17'd53549: data = 8'hca;
      17'd53550: data = 8'hce;
      17'd53551: data = 8'hc9;
      17'd53552: data = 8'hbc;
      17'd53553: data = 8'hc0;
      17'd53554: data = 8'hc6;
      17'd53555: data = 8'hc4;
      17'd53556: data = 8'hc6;
      17'd53557: data = 8'hd8;
      17'd53558: data = 8'hda;
      17'd53559: data = 8'hd6;
      17'd53560: data = 8'hdc;
      17'd53561: data = 8'he2;
      17'd53562: data = 8'hdb;
      17'd53563: data = 8'hda;
      17'd53564: data = 8'he9;
      17'd53565: data = 8'hef;
      17'd53566: data = 8'hef;
      17'd53567: data = 8'hf6;
      17'd53568: data = 8'hf9;
      17'd53569: data = 8'hf5;
      17'd53570: data = 8'hf2;
      17'd53571: data = 8'hf6;
      17'd53572: data = 8'hfd;
      17'd53573: data = 8'hfd;
      17'd53574: data = 8'h04;
      17'd53575: data = 8'h0c;
      17'd53576: data = 8'h0d;
      17'd53577: data = 8'h12;
      17'd53578: data = 8'h12;
      17'd53579: data = 8'h0d;
      17'd53580: data = 8'h0a;
      17'd53581: data = 8'h0e;
      17'd53582: data = 8'h12;
      17'd53583: data = 8'h12;
      17'd53584: data = 8'h15;
      17'd53585: data = 8'h15;
      17'd53586: data = 8'h12;
      17'd53587: data = 8'h0a;
      17'd53588: data = 8'h09;
      17'd53589: data = 8'h0a;
      17'd53590: data = 8'h06;
      17'd53591: data = 8'h06;
      17'd53592: data = 8'h05;
      17'd53593: data = 8'h05;
      17'd53594: data = 8'h02;
      17'd53595: data = 8'hfd;
      17'd53596: data = 8'hfa;
      17'd53597: data = 8'hf9;
      17'd53598: data = 8'hf4;
      17'd53599: data = 8'hf1;
      17'd53600: data = 8'hf6;
      17'd53601: data = 8'hf5;
      17'd53602: data = 8'hf2;
      17'd53603: data = 8'hf1;
      17'd53604: data = 8'hed;
      17'd53605: data = 8'hec;
      17'd53606: data = 8'hed;
      17'd53607: data = 8'hf1;
      17'd53608: data = 8'hf2;
      17'd53609: data = 8'hf1;
      17'd53610: data = 8'hf2;
      17'd53611: data = 8'hf5;
      17'd53612: data = 8'hf2;
      17'd53613: data = 8'hf2;
      17'd53614: data = 8'hf6;
      17'd53615: data = 8'hf6;
      17'd53616: data = 8'hf4;
      17'd53617: data = 8'hfc;
      17'd53618: data = 8'hfe;
      17'd53619: data = 8'hfd;
      17'd53620: data = 8'hfd;
      17'd53621: data = 8'hfe;
      17'd53622: data = 8'hfd;
      17'd53623: data = 8'hfc;
      17'd53624: data = 8'h00;
      17'd53625: data = 8'h05;
      17'd53626: data = 8'h0a;
      17'd53627: data = 8'h0c;
      17'd53628: data = 8'h0e;
      17'd53629: data = 8'h11;
      17'd53630: data = 8'h13;
      17'd53631: data = 8'h12;
      17'd53632: data = 8'h15;
      17'd53633: data = 8'h1b;
      17'd53634: data = 8'h1e;
      17'd53635: data = 8'h22;
      17'd53636: data = 8'h1e;
      17'd53637: data = 8'h1a;
      17'd53638: data = 8'h16;
      17'd53639: data = 8'h15;
      17'd53640: data = 8'h12;
      17'd53641: data = 8'h13;
      17'd53642: data = 8'h1b;
      17'd53643: data = 8'h19;
      17'd53644: data = 8'h15;
      17'd53645: data = 8'h16;
      17'd53646: data = 8'h1a;
      17'd53647: data = 8'h11;
      17'd53648: data = 8'h0c;
      17'd53649: data = 8'h11;
      17'd53650: data = 8'h11;
      17'd53651: data = 8'h12;
      17'd53652: data = 8'h13;
      17'd53653: data = 8'h19;
      17'd53654: data = 8'h13;
      17'd53655: data = 8'h0c;
      17'd53656: data = 8'h0c;
      17'd53657: data = 8'h06;
      17'd53658: data = 8'h04;
      17'd53659: data = 8'h00;
      17'd53660: data = 8'h01;
      17'd53661: data = 8'h06;
      17'd53662: data = 8'h0a;
      17'd53663: data = 8'h09;
      17'd53664: data = 8'h06;
      17'd53665: data = 8'h00;
      17'd53666: data = 8'hf5;
      17'd53667: data = 8'hef;
      17'd53668: data = 8'he7;
      17'd53669: data = 8'he7;
      17'd53670: data = 8'hec;
      17'd53671: data = 8'hf1;
      17'd53672: data = 8'hf5;
      17'd53673: data = 8'hf6;
      17'd53674: data = 8'hfa;
      17'd53675: data = 8'hf4;
      17'd53676: data = 8'hf4;
      17'd53677: data = 8'hfd;
      17'd53678: data = 8'h0a;
      17'd53679: data = 8'h0e;
      17'd53680: data = 8'h1b;
      17'd53681: data = 8'h2d;
      17'd53682: data = 8'h2d;
      17'd53683: data = 8'h2b;
      17'd53684: data = 8'h23;
      17'd53685: data = 8'h1e;
      17'd53686: data = 8'h1a;
      17'd53687: data = 8'h1b;
      17'd53688: data = 8'h22;
      17'd53689: data = 8'h23;
      17'd53690: data = 8'h27;
      17'd53691: data = 8'h23;
      17'd53692: data = 8'h1c;
      17'd53693: data = 8'h1b;
      17'd53694: data = 8'h19;
      17'd53695: data = 8'h16;
      17'd53696: data = 8'h1b;
      17'd53697: data = 8'h26;
      17'd53698: data = 8'h2d;
      17'd53699: data = 8'h31;
      17'd53700: data = 8'h34;
      17'd53701: data = 8'h2d;
      17'd53702: data = 8'h23;
      17'd53703: data = 8'h1c;
      17'd53704: data = 8'h16;
      17'd53705: data = 8'h11;
      17'd53706: data = 8'h0e;
      17'd53707: data = 8'h0c;
      17'd53708: data = 8'h0a;
      17'd53709: data = 8'h02;
      17'd53710: data = 8'hf9;
      17'd53711: data = 8'hed;
      17'd53712: data = 8'he5;
      17'd53713: data = 8'he0;
      17'd53714: data = 8'he0;
      17'd53715: data = 8'he5;
      17'd53716: data = 8'he4;
      17'd53717: data = 8'he5;
      17'd53718: data = 8'he4;
      17'd53719: data = 8'he0;
      17'd53720: data = 8'hda;
      17'd53721: data = 8'hd1;
      17'd53722: data = 8'hd1;
      17'd53723: data = 8'hd1;
      17'd53724: data = 8'hd1;
      17'd53725: data = 8'hd2;
      17'd53726: data = 8'hd3;
      17'd53727: data = 8'hd1;
      17'd53728: data = 8'hcb;
      17'd53729: data = 8'hc6;
      17'd53730: data = 8'hc4;
      17'd53731: data = 8'hc6;
      17'd53732: data = 8'hc9;
      17'd53733: data = 8'hd3;
      17'd53734: data = 8'he0;
      17'd53735: data = 8'he3;
      17'd53736: data = 8'he7;
      17'd53737: data = 8'hec;
      17'd53738: data = 8'hf2;
      17'd53739: data = 8'hf6;
      17'd53740: data = 8'hfe;
      17'd53741: data = 8'h02;
      17'd53742: data = 8'h09;
      17'd53743: data = 8'h0e;
      17'd53744: data = 8'h12;
      17'd53745: data = 8'h12;
      17'd53746: data = 8'h0e;
      17'd53747: data = 8'h11;
      17'd53748: data = 8'h12;
      17'd53749: data = 8'h13;
      17'd53750: data = 8'h19;
      17'd53751: data = 8'h1c;
      17'd53752: data = 8'h22;
      17'd53753: data = 8'h27;
      17'd53754: data = 8'h2b;
      17'd53755: data = 8'h2c;
      17'd53756: data = 8'h2d;
      17'd53757: data = 8'h2f;
      17'd53758: data = 8'h34;
      17'd53759: data = 8'h36;
      17'd53760: data = 8'h39;
      17'd53761: data = 8'h36;
      17'd53762: data = 8'h36;
      17'd53763: data = 8'h31;
      17'd53764: data = 8'h29;
      17'd53765: data = 8'h22;
      17'd53766: data = 8'h1a;
      17'd53767: data = 8'h13;
      17'd53768: data = 8'h12;
      17'd53769: data = 8'h0e;
      17'd53770: data = 8'h0d;
      17'd53771: data = 8'h06;
      17'd53772: data = 8'h01;
      17'd53773: data = 8'hfd;
      17'd53774: data = 8'hf9;
      17'd53775: data = 8'hf6;
      17'd53776: data = 8'hf6;
      17'd53777: data = 8'hf5;
      17'd53778: data = 8'hf4;
      17'd53779: data = 8'hf2;
      17'd53780: data = 8'hec;
      17'd53781: data = 8'he5;
      17'd53782: data = 8'hde;
      17'd53783: data = 8'hda;
      17'd53784: data = 8'hd5;
      17'd53785: data = 8'hce;
      17'd53786: data = 8'hcb;
      17'd53787: data = 8'hcb;
      17'd53788: data = 8'hcb;
      17'd53789: data = 8'hca;
      17'd53790: data = 8'hca;
      17'd53791: data = 8'hc9;
      17'd53792: data = 8'hcb;
      17'd53793: data = 8'hc9;
      17'd53794: data = 8'hc6;
      17'd53795: data = 8'hce;
      17'd53796: data = 8'hd1;
      17'd53797: data = 8'hcd;
      17'd53798: data = 8'hd3;
      17'd53799: data = 8'hd6;
      17'd53800: data = 8'hd2;
      17'd53801: data = 8'hd3;
      17'd53802: data = 8'hd8;
      17'd53803: data = 8'hda;
      17'd53804: data = 8'hd5;
      17'd53805: data = 8'hd8;
      17'd53806: data = 8'he0;
      17'd53807: data = 8'he0;
      17'd53808: data = 8'he3;
      17'd53809: data = 8'he9;
      17'd53810: data = 8'heb;
      17'd53811: data = 8'heb;
      17'd53812: data = 8'hed;
      17'd53813: data = 8'hf4;
      17'd53814: data = 8'hf4;
      17'd53815: data = 8'hf5;
      17'd53816: data = 8'hfa;
      17'd53817: data = 8'hfe;
      17'd53818: data = 8'hfe;
      17'd53819: data = 8'h01;
      17'd53820: data = 8'h05;
      17'd53821: data = 8'h05;
      17'd53822: data = 8'h04;
      17'd53823: data = 8'h05;
      17'd53824: data = 8'h0a;
      17'd53825: data = 8'h09;
      17'd53826: data = 8'h09;
      17'd53827: data = 8'h0c;
      17'd53828: data = 8'h0c;
      17'd53829: data = 8'h0d;
      17'd53830: data = 8'h0d;
      17'd53831: data = 8'h0c;
      17'd53832: data = 8'h0a;
      17'd53833: data = 8'h09;
      17'd53834: data = 8'h09;
      17'd53835: data = 8'h0a;
      17'd53836: data = 8'h09;
      17'd53837: data = 8'h0a;
      17'd53838: data = 8'h0a;
      17'd53839: data = 8'h09;
      17'd53840: data = 8'h04;
      17'd53841: data = 8'h02;
      17'd53842: data = 8'h01;
      17'd53843: data = 8'h00;
      17'd53844: data = 8'h00;
      17'd53845: data = 8'h02;
      17'd53846: data = 8'h02;
      17'd53847: data = 8'h01;
      17'd53848: data = 8'h01;
      17'd53849: data = 8'h01;
      17'd53850: data = 8'hfd;
      17'd53851: data = 8'hfc;
      17'd53852: data = 8'h00;
      17'd53853: data = 8'h00;
      17'd53854: data = 8'hfd;
      17'd53855: data = 8'h00;
      17'd53856: data = 8'h00;
      17'd53857: data = 8'hfa;
      17'd53858: data = 8'hf9;
      17'd53859: data = 8'hfc;
      17'd53860: data = 8'hfc;
      17'd53861: data = 8'hf6;
      17'd53862: data = 8'hfa;
      17'd53863: data = 8'hfd;
      17'd53864: data = 8'hfc;
      17'd53865: data = 8'hfd;
      17'd53866: data = 8'h00;
      17'd53867: data = 8'h02;
      17'd53868: data = 8'h02;
      17'd53869: data = 8'h05;
      17'd53870: data = 8'h0a;
      17'd53871: data = 8'h0a;
      17'd53872: data = 8'h0a;
      17'd53873: data = 8'h0a;
      17'd53874: data = 8'h0a;
      17'd53875: data = 8'h09;
      17'd53876: data = 8'h09;
      17'd53877: data = 8'h09;
      17'd53878: data = 8'h05;
      17'd53879: data = 8'h0c;
      17'd53880: data = 8'h0d;
      17'd53881: data = 8'h0e;
      17'd53882: data = 8'h0a;
      17'd53883: data = 8'h0d;
      17'd53884: data = 8'h0e;
      17'd53885: data = 8'h0d;
      17'd53886: data = 8'h0e;
      17'd53887: data = 8'h16;
      17'd53888: data = 8'h19;
      17'd53889: data = 8'h13;
      17'd53890: data = 8'h15;
      17'd53891: data = 8'h16;
      17'd53892: data = 8'h13;
      17'd53893: data = 8'h0a;
      17'd53894: data = 8'h0d;
      17'd53895: data = 8'h13;
      17'd53896: data = 8'h11;
      17'd53897: data = 8'h11;
      17'd53898: data = 8'h13;
      17'd53899: data = 8'h12;
      17'd53900: data = 8'h06;
      17'd53901: data = 8'h09;
      17'd53902: data = 8'h09;
      17'd53903: data = 8'h04;
      17'd53904: data = 8'h09;
      17'd53905: data = 8'h09;
      17'd53906: data = 8'h00;
      17'd53907: data = 8'hfc;
      17'd53908: data = 8'hfc;
      17'd53909: data = 8'hf9;
      17'd53910: data = 8'hef;
      17'd53911: data = 8'hf4;
      17'd53912: data = 8'hfd;
      17'd53913: data = 8'hf9;
      17'd53914: data = 8'hf6;
      17'd53915: data = 8'h01;
      17'd53916: data = 8'h02;
      17'd53917: data = 8'hfe;
      17'd53918: data = 8'h04;
      17'd53919: data = 8'h0e;
      17'd53920: data = 8'h12;
      17'd53921: data = 8'h16;
      17'd53922: data = 8'h1a;
      17'd53923: data = 8'h1b;
      17'd53924: data = 8'h19;
      17'd53925: data = 8'h12;
      17'd53926: data = 8'h0e;
      17'd53927: data = 8'h0d;
      17'd53928: data = 8'h09;
      17'd53929: data = 8'h0c;
      17'd53930: data = 8'h11;
      17'd53931: data = 8'h13;
      17'd53932: data = 8'h11;
      17'd53933: data = 8'h15;
      17'd53934: data = 8'h15;
      17'd53935: data = 8'h11;
      17'd53936: data = 8'h16;
      17'd53937: data = 8'h24;
      17'd53938: data = 8'h27;
      17'd53939: data = 8'h27;
      17'd53940: data = 8'h2c;
      17'd53941: data = 8'h2b;
      17'd53942: data = 8'h22;
      17'd53943: data = 8'h19;
      17'd53944: data = 8'h16;
      17'd53945: data = 8'h11;
      17'd53946: data = 8'h0a;
      17'd53947: data = 8'h0a;
      17'd53948: data = 8'h0c;
      17'd53949: data = 8'h0a;
      17'd53950: data = 8'h02;
      17'd53951: data = 8'hfe;
      17'd53952: data = 8'hfe;
      17'd53953: data = 8'hf6;
      17'd53954: data = 8'hf1;
      17'd53955: data = 8'hf5;
      17'd53956: data = 8'hf9;
      17'd53957: data = 8'hf4;
      17'd53958: data = 8'hf2;
      17'd53959: data = 8'hf1;
      17'd53960: data = 8'he5;
      17'd53961: data = 8'hdc;
      17'd53962: data = 8'hda;
      17'd53963: data = 8'hd5;
      17'd53964: data = 8'hd3;
      17'd53965: data = 8'hd3;
      17'd53966: data = 8'hd5;
      17'd53967: data = 8'hd3;
      17'd53968: data = 8'hd1;
      17'd53969: data = 8'hcb;
      17'd53970: data = 8'hca;
      17'd53971: data = 8'hcd;
      17'd53972: data = 8'hd1;
      17'd53973: data = 8'hd5;
      17'd53974: data = 8'he0;
      17'd53975: data = 8'he4;
      17'd53976: data = 8'he9;
      17'd53977: data = 8'hef;
      17'd53978: data = 8'hef;
      17'd53979: data = 8'hed;
      17'd53980: data = 8'hef;
      17'd53981: data = 8'hf4;
      17'd53982: data = 8'hf4;
      17'd53983: data = 8'hf9;
      17'd53984: data = 8'hfe;
      17'd53985: data = 8'h00;
      17'd53986: data = 8'hfd;
      17'd53987: data = 8'hfe;
      17'd53988: data = 8'h04;
      17'd53989: data = 8'h06;
      17'd53990: data = 8'h0c;
      17'd53991: data = 8'h13;
      17'd53992: data = 8'h1c;
      17'd53993: data = 8'h22;
      17'd53994: data = 8'h24;
      17'd53995: data = 8'h24;
      17'd53996: data = 8'h26;
      17'd53997: data = 8'h26;
      17'd53998: data = 8'h24;
      17'd53999: data = 8'h27;
      17'd54000: data = 8'h26;
      17'd54001: data = 8'h24;
      17'd54002: data = 8'h24;
      17'd54003: data = 8'h1f;
      17'd54004: data = 8'h1b;
      17'd54005: data = 8'h19;
      17'd54006: data = 8'h19;
      17'd54007: data = 8'h16;
      17'd54008: data = 8'h16;
      17'd54009: data = 8'h16;
      17'd54010: data = 8'h16;
      17'd54011: data = 8'h15;
      17'd54012: data = 8'h0e;
      17'd54013: data = 8'h0c;
      17'd54014: data = 8'h0a;
      17'd54015: data = 8'h06;
      17'd54016: data = 8'h04;
      17'd54017: data = 8'h00;
      17'd54018: data = 8'hf9;
      17'd54019: data = 8'hf4;
      17'd54020: data = 8'hf1;
      17'd54021: data = 8'hec;
      17'd54022: data = 8'he4;
      17'd54023: data = 8'he3;
      17'd54024: data = 8'he9;
      17'd54025: data = 8'he5;
      17'd54026: data = 8'he0;
      17'd54027: data = 8'hde;
      17'd54028: data = 8'he2;
      17'd54029: data = 8'hde;
      17'd54030: data = 8'hd5;
      17'd54031: data = 8'hd2;
      17'd54032: data = 8'hdc;
      17'd54033: data = 8'he0;
      17'd54034: data = 8'hd5;
      17'd54035: data = 8'hd6;
      17'd54036: data = 8'he0;
      17'd54037: data = 8'hd6;
      17'd54038: data = 8'hc6;
      17'd54039: data = 8'hcd;
      17'd54040: data = 8'hd3;
      17'd54041: data = 8'hcd;
      17'd54042: data = 8'hd2;
      17'd54043: data = 8'hdc;
      17'd54044: data = 8'hd6;
      17'd54045: data = 8'hd1;
      17'd54046: data = 8'hdb;
      17'd54047: data = 8'hdb;
      17'd54048: data = 8'hd3;
      17'd54049: data = 8'hdc;
      17'd54050: data = 8'hed;
      17'd54051: data = 8'he7;
      17'd54052: data = 8'he3;
      17'd54053: data = 8'hef;
      17'd54054: data = 8'hf5;
      17'd54055: data = 8'heb;
      17'd54056: data = 8'he7;
      17'd54057: data = 8'hed;
      17'd54058: data = 8'hec;
      17'd54059: data = 8'hec;
      17'd54060: data = 8'hf5;
      17'd54061: data = 8'h00;
      17'd54062: data = 8'h01;
      17'd54063: data = 8'h00;
      17'd54064: data = 8'h02;
      17'd54065: data = 8'h01;
      17'd54066: data = 8'hfe;
      17'd54067: data = 8'h02;
      17'd54068: data = 8'h06;
      17'd54069: data = 8'h09;
      17'd54070: data = 8'h06;
      17'd54071: data = 8'h0a;
      17'd54072: data = 8'h0a;
      17'd54073: data = 8'h02;
      17'd54074: data = 8'hfd;
      17'd54075: data = 8'hfe;
      17'd54076: data = 8'h02;
      17'd54077: data = 8'h02;
      17'd54078: data = 8'h06;
      17'd54079: data = 8'h0c;
      17'd54080: data = 8'h0d;
      17'd54081: data = 8'h0a;
      17'd54082: data = 8'h05;
      17'd54083: data = 8'h06;
      17'd54084: data = 8'h05;
      17'd54085: data = 8'h05;
      17'd54086: data = 8'h06;
      17'd54087: data = 8'h06;
      17'd54088: data = 8'h05;
      17'd54089: data = 8'h05;
      17'd54090: data = 8'h05;
      17'd54091: data = 8'h00;
      17'd54092: data = 8'h00;
      17'd54093: data = 8'h04;
      17'd54094: data = 8'h05;
      17'd54095: data = 8'h05;
      17'd54096: data = 8'h06;
      17'd54097: data = 8'h0a;
      17'd54098: data = 8'h0a;
      17'd54099: data = 8'h05;
      17'd54100: data = 8'h04;
      17'd54101: data = 8'h06;
      17'd54102: data = 8'h09;
      17'd54103: data = 8'h02;
      17'd54104: data = 8'h06;
      17'd54105: data = 8'h11;
      17'd54106: data = 8'h0c;
      17'd54107: data = 8'h06;
      17'd54108: data = 8'h05;
      17'd54109: data = 8'h09;
      17'd54110: data = 8'h06;
      17'd54111: data = 8'h05;
      17'd54112: data = 8'h04;
      17'd54113: data = 8'h09;
      17'd54114: data = 8'h0a;
      17'd54115: data = 8'h0c;
      17'd54116: data = 8'h06;
      17'd54117: data = 8'h05;
      17'd54118: data = 8'h09;
      17'd54119: data = 8'h05;
      17'd54120: data = 8'h09;
      17'd54121: data = 8'h0d;
      17'd54122: data = 8'h0e;
      17'd54123: data = 8'h09;
      17'd54124: data = 8'h11;
      17'd54125: data = 8'h0e;
      17'd54126: data = 8'h09;
      17'd54127: data = 8'h05;
      17'd54128: data = 8'h0a;
      17'd54129: data = 8'h09;
      17'd54130: data = 8'h05;
      17'd54131: data = 8'h09;
      17'd54132: data = 8'h11;
      17'd54133: data = 8'h0c;
      17'd54134: data = 8'h05;
      17'd54135: data = 8'h12;
      17'd54136: data = 8'h0c;
      17'd54137: data = 8'h00;
      17'd54138: data = 8'h0a;
      17'd54139: data = 8'h19;
      17'd54140: data = 8'h11;
      17'd54141: data = 8'h0e;
      17'd54142: data = 8'h13;
      17'd54143: data = 8'h0a;
      17'd54144: data = 8'hf9;
      17'd54145: data = 8'hf4;
      17'd54146: data = 8'hf5;
      17'd54147: data = 8'hf2;
      17'd54148: data = 8'hf6;
      17'd54149: data = 8'h00;
      17'd54150: data = 8'h05;
      17'd54151: data = 8'h02;
      17'd54152: data = 8'h02;
      17'd54153: data = 8'h04;
      17'd54154: data = 8'h01;
      17'd54155: data = 8'hfe;
      17'd54156: data = 8'h0a;
      17'd54157: data = 8'h19;
      17'd54158: data = 8'h1b;
      17'd54159: data = 8'h19;
      17'd54160: data = 8'h19;
      17'd54161: data = 8'h16;
      17'd54162: data = 8'h09;
      17'd54163: data = 8'h00;
      17'd54164: data = 8'h06;
      17'd54165: data = 8'h09;
      17'd54166: data = 8'h06;
      17'd54167: data = 8'h12;
      17'd54168: data = 8'h19;
      17'd54169: data = 8'h16;
      17'd54170: data = 8'h1a;
      17'd54171: data = 8'h1b;
      17'd54172: data = 8'h12;
      17'd54173: data = 8'h15;
      17'd54174: data = 8'h1e;
      17'd54175: data = 8'h22;
      17'd54176: data = 8'h23;
      17'd54177: data = 8'h29;
      17'd54178: data = 8'h29;
      17'd54179: data = 8'h23;
      17'd54180: data = 8'h1b;
      17'd54181: data = 8'h12;
      17'd54182: data = 8'h0e;
      17'd54183: data = 8'h0d;
      17'd54184: data = 8'h0c;
      17'd54185: data = 8'h09;
      17'd54186: data = 8'h0d;
      17'd54187: data = 8'h13;
      17'd54188: data = 8'h06;
      17'd54189: data = 8'h00;
      17'd54190: data = 8'h04;
      17'd54191: data = 8'h01;
      17'd54192: data = 8'hfc;
      17'd54193: data = 8'hfd;
      17'd54194: data = 8'h00;
      17'd54195: data = 8'hfe;
      17'd54196: data = 8'hfc;
      17'd54197: data = 8'hf4;
      17'd54198: data = 8'hef;
      17'd54199: data = 8'he7;
      17'd54200: data = 8'hdc;
      17'd54201: data = 8'hdb;
      17'd54202: data = 8'hd8;
      17'd54203: data = 8'hd5;
      17'd54204: data = 8'hd6;
      17'd54205: data = 8'hdb;
      17'd54206: data = 8'hd8;
      17'd54207: data = 8'hd5;
      17'd54208: data = 8'hdb;
      17'd54209: data = 8'he0;
      17'd54210: data = 8'he0;
      17'd54211: data = 8'he4;
      17'd54212: data = 8'he9;
      17'd54213: data = 8'heb;
      17'd54214: data = 8'he9;
      17'd54215: data = 8'he9;
      17'd54216: data = 8'he9;
      17'd54217: data = 8'he4;
      17'd54218: data = 8'he7;
      17'd54219: data = 8'he9;
      17'd54220: data = 8'he7;
      17'd54221: data = 8'hed;
      17'd54222: data = 8'hf2;
      17'd54223: data = 8'hf4;
      17'd54224: data = 8'hfa;
      17'd54225: data = 8'hfd;
      17'd54226: data = 8'h01;
      17'd54227: data = 8'h06;
      17'd54228: data = 8'h0d;
      17'd54229: data = 8'h11;
      17'd54230: data = 8'h13;
      17'd54231: data = 8'h16;
      17'd54232: data = 8'h19;
      17'd54233: data = 8'h15;
      17'd54234: data = 8'h13;
      17'd54235: data = 8'h15;
      17'd54236: data = 8'h13;
      17'd54237: data = 8'h13;
      17'd54238: data = 8'h1a;
      17'd54239: data = 8'h1b;
      17'd54240: data = 8'h1a;
      17'd54241: data = 8'h1c;
      17'd54242: data = 8'h1b;
      17'd54243: data = 8'h1a;
      17'd54244: data = 8'h1a;
      17'd54245: data = 8'h19;
      17'd54246: data = 8'h1a;
      17'd54247: data = 8'h1e;
      17'd54248: data = 8'h1c;
      17'd54249: data = 8'h1a;
      17'd54250: data = 8'h15;
      17'd54251: data = 8'h0e;
      17'd54252: data = 8'h0d;
      17'd54253: data = 8'h09;
      17'd54254: data = 8'h05;
      17'd54255: data = 8'h02;
      17'd54256: data = 8'h04;
      17'd54257: data = 8'h05;
      17'd54258: data = 8'h04;
      17'd54259: data = 8'h01;
      17'd54260: data = 8'hfe;
      17'd54261: data = 8'hfc;
      17'd54262: data = 8'hf4;
      17'd54263: data = 8'hef;
      17'd54264: data = 8'hed;
      17'd54265: data = 8'hef;
      17'd54266: data = 8'hed;
      17'd54267: data = 8'hec;
      17'd54268: data = 8'he9;
      17'd54269: data = 8'heb;
      17'd54270: data = 8'he7;
      17'd54271: data = 8'he0;
      17'd54272: data = 8'hdb;
      17'd54273: data = 8'hdb;
      17'd54274: data = 8'hdb;
      17'd54275: data = 8'hda;
      17'd54276: data = 8'hda;
      17'd54277: data = 8'hdb;
      17'd54278: data = 8'hdc;
      17'd54279: data = 8'hd8;
      17'd54280: data = 8'hd6;
      17'd54281: data = 8'hd6;
      17'd54282: data = 8'hd3;
      17'd54283: data = 8'hd5;
      17'd54284: data = 8'hda;
      17'd54285: data = 8'hd6;
      17'd54286: data = 8'hd8;
      17'd54287: data = 8'he0;
      17'd54288: data = 8'hde;
      17'd54289: data = 8'hd8;
      17'd54290: data = 8'hd8;
      17'd54291: data = 8'he0;
      17'd54292: data = 8'hda;
      17'd54293: data = 8'hd5;
      17'd54294: data = 8'he2;
      17'd54295: data = 8'he7;
      17'd54296: data = 8'he3;
      17'd54297: data = 8'he5;
      17'd54298: data = 8'hef;
      17'd54299: data = 8'hef;
      17'd54300: data = 8'hf1;
      17'd54301: data = 8'hf4;
      17'd54302: data = 8'hf4;
      17'd54303: data = 8'hf5;
      17'd54304: data = 8'hf6;
      17'd54305: data = 8'hfc;
      17'd54306: data = 8'hf9;
      17'd54307: data = 8'hf6;
      17'd54308: data = 8'hf6;
      17'd54309: data = 8'hf5;
      17'd54310: data = 8'hf5;
      17'd54311: data = 8'hf6;
      17'd54312: data = 8'hfa;
      17'd54313: data = 8'hfc;
      17'd54314: data = 8'hfd;
      17'd54315: data = 8'hfe;
      17'd54316: data = 8'h01;
      17'd54317: data = 8'h05;
      17'd54318: data = 8'h02;
      17'd54319: data = 8'h01;
      17'd54320: data = 8'h04;
      17'd54321: data = 8'h05;
      17'd54322: data = 8'h05;
      17'd54323: data = 8'h05;
      17'd54324: data = 8'h06;
      17'd54325: data = 8'h0a;
      17'd54326: data = 8'h09;
      17'd54327: data = 8'h0a;
      17'd54328: data = 8'h0c;
      17'd54329: data = 8'h0a;
      17'd54330: data = 8'h09;
      17'd54331: data = 8'h0a;
      17'd54332: data = 8'h0c;
      17'd54333: data = 8'h0c;
      17'd54334: data = 8'h0c;
      17'd54335: data = 8'h0d;
      17'd54336: data = 8'h0e;
      17'd54337: data = 8'h09;
      17'd54338: data = 8'h0c;
      17'd54339: data = 8'h11;
      17'd54340: data = 8'h0e;
      17'd54341: data = 8'h0d;
      17'd54342: data = 8'h12;
      17'd54343: data = 8'h13;
      17'd54344: data = 8'h0d;
      17'd54345: data = 8'h11;
      17'd54346: data = 8'h16;
      17'd54347: data = 8'h0e;
      17'd54348: data = 8'h0a;
      17'd54349: data = 8'h0e;
      17'd54350: data = 8'h13;
      17'd54351: data = 8'h0a;
      17'd54352: data = 8'h0a;
      17'd54353: data = 8'h0c;
      17'd54354: data = 8'h06;
      17'd54355: data = 8'h00;
      17'd54356: data = 8'h05;
      17'd54357: data = 8'h0e;
      17'd54358: data = 8'h02;
      17'd54359: data = 8'h01;
      17'd54360: data = 8'h0d;
      17'd54361: data = 8'h09;
      17'd54362: data = 8'h04;
      17'd54363: data = 8'h02;
      17'd54364: data = 8'h05;
      17'd54365: data = 8'h05;
      17'd54366: data = 8'h04;
      17'd54367: data = 8'h0a;
      17'd54368: data = 8'h02;
      17'd54369: data = 8'h02;
      17'd54370: data = 8'h04;
      17'd54371: data = 8'h01;
      17'd54372: data = 8'hfd;
      17'd54373: data = 8'h04;
      17'd54374: data = 8'h06;
      17'd54375: data = 8'h06;
      17'd54376: data = 8'h0a;
      17'd54377: data = 8'h0c;
      17'd54378: data = 8'h0a;
      17'd54379: data = 8'h06;
      17'd54380: data = 8'h04;
      17'd54381: data = 8'h01;
      17'd54382: data = 8'hfe;
      17'd54383: data = 8'hfa;
      17'd54384: data = 8'hf9;
      17'd54385: data = 8'hef;
      17'd54386: data = 8'hf4;
      17'd54387: data = 8'hfa;
      17'd54388: data = 8'hfc;
      17'd54389: data = 8'hfe;
      17'd54390: data = 8'h09;
      17'd54391: data = 8'h06;
      17'd54392: data = 8'h0d;
      17'd54393: data = 8'h11;
      17'd54394: data = 8'h0c;
      17'd54395: data = 8'h11;
      17'd54396: data = 8'h0e;
      17'd54397: data = 8'h0e;
      17'd54398: data = 8'h13;
      17'd54399: data = 8'h11;
      17'd54400: data = 8'h0e;
      17'd54401: data = 8'h13;
      17'd54402: data = 8'h09;
      17'd54403: data = 8'h02;
      17'd54404: data = 8'h0a;
      17'd54405: data = 8'h09;
      17'd54406: data = 8'h0c;
      17'd54407: data = 8'h12;
      17'd54408: data = 8'h15;
      17'd54409: data = 8'h22;
      17'd54410: data = 8'h1f;
      17'd54411: data = 8'h1a;
      17'd54412: data = 8'h1f;
      17'd54413: data = 8'h1b;
      17'd54414: data = 8'h15;
      17'd54415: data = 8'h1c;
      17'd54416: data = 8'h1b;
      17'd54417: data = 8'h19;
      17'd54418: data = 8'h1e;
      17'd54419: data = 8'h1c;
      17'd54420: data = 8'h12;
      17'd54421: data = 8'h0c;
      17'd54422: data = 8'h0a;
      17'd54423: data = 8'h0d;
      17'd54424: data = 8'h06;
      17'd54425: data = 8'h02;
      17'd54426: data = 8'h12;
      17'd54427: data = 8'h0e;
      17'd54428: data = 8'h0c;
      17'd54429: data = 8'h0d;
      17'd54430: data = 8'h06;
      17'd54431: data = 8'h00;
      17'd54432: data = 8'hfe;
      17'd54433: data = 8'hfa;
      17'd54434: data = 8'hf6;
      17'd54435: data = 8'hf9;
      17'd54436: data = 8'hf5;
      17'd54437: data = 8'hf5;
      17'd54438: data = 8'hf1;
      17'd54439: data = 8'he7;
      17'd54440: data = 8'he5;
      17'd54441: data = 8'he2;
      17'd54442: data = 8'hdb;
      17'd54443: data = 8'hde;
      17'd54444: data = 8'he3;
      17'd54445: data = 8'he4;
      17'd54446: data = 8'he7;
      17'd54447: data = 8'he7;
      17'd54448: data = 8'he7;
      17'd54449: data = 8'he4;
      17'd54450: data = 8'he0;
      17'd54451: data = 8'he0;
      17'd54452: data = 8'he3;
      17'd54453: data = 8'he4;
      17'd54454: data = 8'he5;
      17'd54455: data = 8'he9;
      17'd54456: data = 8'he9;
      17'd54457: data = 8'he9;
      17'd54458: data = 8'heb;
      17'd54459: data = 8'he5;
      17'd54460: data = 8'he9;
      17'd54461: data = 8'hf1;
      17'd54462: data = 8'hf2;
      17'd54463: data = 8'hf9;
      17'd54464: data = 8'hfd;
      17'd54465: data = 8'hfe;
      17'd54466: data = 8'h01;
      17'd54467: data = 8'h04;
      17'd54468: data = 8'h01;
      17'd54469: data = 8'h02;
      17'd54470: data = 8'h05;
      17'd54471: data = 8'h04;
      17'd54472: data = 8'h09;
      17'd54473: data = 8'h0a;
      17'd54474: data = 8'h0a;
      17'd54475: data = 8'h0d;
      17'd54476: data = 8'h0d;
      17'd54477: data = 8'h0a;
      17'd54478: data = 8'h0d;
      17'd54479: data = 8'h12;
      17'd54480: data = 8'h19;
      17'd54481: data = 8'h19;
      17'd54482: data = 8'h1b;
      17'd54483: data = 8'h1e;
      17'd54484: data = 8'h1b;
      17'd54485: data = 8'h1a;
      17'd54486: data = 8'h16;
      17'd54487: data = 8'h13;
      17'd54488: data = 8'h11;
      17'd54489: data = 8'h11;
      17'd54490: data = 8'h0d;
      17'd54491: data = 8'h0d;
      17'd54492: data = 8'h0d;
      17'd54493: data = 8'h0d;
      17'd54494: data = 8'h0c;
      17'd54495: data = 8'h06;
      17'd54496: data = 8'h05;
      17'd54497: data = 8'h0a;
      17'd54498: data = 8'h06;
      17'd54499: data = 8'h06;
      17'd54500: data = 8'h06;
      17'd54501: data = 8'h05;
      17'd54502: data = 8'h04;
      17'd54503: data = 8'h01;
      17'd54504: data = 8'hf6;
      17'd54505: data = 8'hed;
      17'd54506: data = 8'hf1;
      17'd54507: data = 8'hed;
      17'd54508: data = 8'hed;
      17'd54509: data = 8'hed;
      17'd54510: data = 8'hef;
      17'd54511: data = 8'hf5;
      17'd54512: data = 8'hf4;
      17'd54513: data = 8'hed;
      17'd54514: data = 8'hec;
      17'd54515: data = 8'hec;
      17'd54516: data = 8'he9;
      17'd54517: data = 8'he3;
      17'd54518: data = 8'he0;
      17'd54519: data = 8'hec;
      17'd54520: data = 8'he9;
      17'd54521: data = 8'hda;
      17'd54522: data = 8'hdc;
      17'd54523: data = 8'hdc;
      17'd54524: data = 8'hd6;
      17'd54525: data = 8'hd6;
      17'd54526: data = 8'hda;
      17'd54527: data = 8'hdb;
      17'd54528: data = 8'hde;
      17'd54529: data = 8'he5;
      17'd54530: data = 8'he9;
      17'd54531: data = 8'he0;
      17'd54532: data = 8'he0;
      17'd54533: data = 8'he4;
      17'd54534: data = 8'hdc;
      17'd54535: data = 8'hd1;
      17'd54536: data = 8'hdb;
      17'd54537: data = 8'he7;
      17'd54538: data = 8'he2;
      17'd54539: data = 8'he3;
      17'd54540: data = 8'heb;
      17'd54541: data = 8'hef;
      17'd54542: data = 8'heb;
      17'd54543: data = 8'he7;
      17'd54544: data = 8'heb;
      17'd54545: data = 8'hec;
      17'd54546: data = 8'hec;
      17'd54547: data = 8'hf1;
      17'd54548: data = 8'hf2;
      17'd54549: data = 8'hed;
      17'd54550: data = 8'hef;
      17'd54551: data = 8'hef;
      17'd54552: data = 8'heb;
      17'd54553: data = 8'heb;
      17'd54554: data = 8'hef;
      17'd54555: data = 8'hf2;
      17'd54556: data = 8'hf6;
      17'd54557: data = 8'hf2;
      17'd54558: data = 8'hfd;
      17'd54559: data = 8'h04;
      17'd54560: data = 8'hfe;
      17'd54561: data = 8'hfe;
      17'd54562: data = 8'h01;
      17'd54563: data = 8'h04;
      17'd54564: data = 8'h04;
      17'd54565: data = 8'h02;
      17'd54566: data = 8'h05;
      17'd54567: data = 8'h0c;
      17'd54568: data = 8'h0c;
      17'd54569: data = 8'h0a;
      17'd54570: data = 8'h11;
      17'd54571: data = 8'h13;
      17'd54572: data = 8'h12;
      17'd54573: data = 8'h19;
      17'd54574: data = 8'h19;
      17'd54575: data = 8'h19;
      17'd54576: data = 8'h19;
      17'd54577: data = 8'h1a;
      17'd54578: data = 8'h15;
      17'd54579: data = 8'h12;
      17'd54580: data = 8'h1b;
      17'd54581: data = 8'h19;
      17'd54582: data = 8'h1b;
      17'd54583: data = 8'h1a;
      17'd54584: data = 8'h16;
      17'd54585: data = 8'h1a;
      17'd54586: data = 8'h16;
      17'd54587: data = 8'h1a;
      17'd54588: data = 8'h1a;
      17'd54589: data = 8'h1b;
      17'd54590: data = 8'h1f;
      17'd54591: data = 8'h1b;
      17'd54592: data = 8'h1f;
      17'd54593: data = 8'h16;
      17'd54594: data = 8'h0c;
      17'd54595: data = 8'h11;
      17'd54596: data = 8'h0a;
      17'd54597: data = 8'h05;
      17'd54598: data = 8'h06;
      17'd54599: data = 8'h0d;
      17'd54600: data = 8'h09;
      17'd54601: data = 8'h06;
      17'd54602: data = 8'h0a;
      17'd54603: data = 8'h05;
      17'd54604: data = 8'h01;
      17'd54605: data = 8'h01;
      17'd54606: data = 8'h05;
      17'd54607: data = 8'h04;
      17'd54608: data = 8'h01;
      17'd54609: data = 8'h0c;
      17'd54610: data = 8'h04;
      17'd54611: data = 8'hfd;
      17'd54612: data = 8'h04;
      17'd54613: data = 8'h00;
      17'd54614: data = 8'hf9;
      17'd54615: data = 8'hfa;
      17'd54616: data = 8'h02;
      17'd54617: data = 8'h06;
      17'd54618: data = 8'h04;
      17'd54619: data = 8'h0d;
      17'd54620: data = 8'h11;
      17'd54621: data = 8'h00;
      17'd54622: data = 8'hfd;
      17'd54623: data = 8'hfd;
      17'd54624: data = 8'hf1;
      17'd54625: data = 8'hed;
      17'd54626: data = 8'hf2;
      17'd54627: data = 8'hf9;
      17'd54628: data = 8'hfa;
      17'd54629: data = 8'hfd;
      17'd54630: data = 8'h01;
      17'd54631: data = 8'h04;
      17'd54632: data = 8'h00;
      17'd54633: data = 8'h00;
      17'd54634: data = 8'h09;
      17'd54635: data = 8'h0d;
      17'd54636: data = 8'h0d;
      17'd54637: data = 8'h15;
      17'd54638: data = 8'h1b;
      17'd54639: data = 8'h1a;
      17'd54640: data = 8'h13;
      17'd54641: data = 8'h0e;
      17'd54642: data = 8'h09;
      17'd54643: data = 8'h02;
      17'd54644: data = 8'h01;
      17'd54645: data = 8'h04;
      17'd54646: data = 8'h0a;
      17'd54647: data = 8'h0e;
      17'd54648: data = 8'h1a;
      17'd54649: data = 8'h1c;
      17'd54650: data = 8'h1a;
      17'd54651: data = 8'h16;
      17'd54652: data = 8'h19;
      17'd54653: data = 8'h1a;
      17'd54654: data = 8'h16;
      17'd54655: data = 8'h1a;
      17'd54656: data = 8'h1f;
      17'd54657: data = 8'h23;
      17'd54658: data = 8'h22;
      17'd54659: data = 8'h1b;
      17'd54660: data = 8'h16;
      17'd54661: data = 8'h0e;
      17'd54662: data = 8'h0a;
      17'd54663: data = 8'h06;
      17'd54664: data = 8'h06;
      17'd54665: data = 8'h0a;
      17'd54666: data = 8'h0c;
      17'd54667: data = 8'h13;
      17'd54668: data = 8'h13;
      17'd54669: data = 8'h0d;
      17'd54670: data = 8'h0a;
      17'd54671: data = 8'h05;
      17'd54672: data = 8'hfe;
      17'd54673: data = 8'hfd;
      17'd54674: data = 8'hfd;
      17'd54675: data = 8'hfd;
      17'd54676: data = 8'hf9;
      17'd54677: data = 8'hf6;
      17'd54678: data = 8'hf5;
      17'd54679: data = 8'hec;
      17'd54680: data = 8'he5;
      17'd54681: data = 8'he2;
      17'd54682: data = 8'hde;
      17'd54683: data = 8'he3;
      17'd54684: data = 8'he9;
      17'd54685: data = 8'hec;
      17'd54686: data = 8'hf1;
      17'd54687: data = 8'hf1;
      17'd54688: data = 8'hed;
      17'd54689: data = 8'hec;
      17'd54690: data = 8'he9;
      17'd54691: data = 8'he4;
      17'd54692: data = 8'he7;
      17'd54693: data = 8'he9;
      17'd54694: data = 8'he9;
      17'd54695: data = 8'heb;
      17'd54696: data = 8'he9;
      17'd54697: data = 8'he9;
      17'd54698: data = 8'he7;
      17'd54699: data = 8'he7;
      17'd54700: data = 8'he9;
      17'd54701: data = 8'hed;
      17'd54702: data = 8'hf4;
      17'd54703: data = 8'hfa;
      17'd54704: data = 8'h00;
      17'd54705: data = 8'h00;
      17'd54706: data = 8'h01;
      17'd54707: data = 8'h00;
      17'd54708: data = 8'hfa;
      17'd54709: data = 8'hfa;
      17'd54710: data = 8'hfa;
      17'd54711: data = 8'hfc;
      17'd54712: data = 8'hfe;
      17'd54713: data = 8'h02;
      17'd54714: data = 8'h04;
      17'd54715: data = 8'h06;
      17'd54716: data = 8'h09;
      17'd54717: data = 8'h06;
      17'd54718: data = 8'h0c;
      17'd54719: data = 8'h0e;
      17'd54720: data = 8'h12;
      17'd54721: data = 8'h19;
      17'd54722: data = 8'h19;
      17'd54723: data = 8'h16;
      17'd54724: data = 8'h15;
      17'd54725: data = 8'h11;
      17'd54726: data = 8'h0c;
      17'd54727: data = 8'h09;
      17'd54728: data = 8'h06;
      17'd54729: data = 8'h0a;
      17'd54730: data = 8'h0a;
      17'd54731: data = 8'h0d;
      17'd54732: data = 8'h0e;
      17'd54733: data = 8'h0d;
      17'd54734: data = 8'h0c;
      17'd54735: data = 8'h0d;
      17'd54736: data = 8'h0c;
      17'd54737: data = 8'h0d;
      17'd54738: data = 8'h0d;
      17'd54739: data = 8'h0e;
      17'd54740: data = 8'h11;
      17'd54741: data = 8'h0d;
      17'd54742: data = 8'h0a;
      17'd54743: data = 8'hfd;
      17'd54744: data = 8'hf1;
      17'd54745: data = 8'heb;
      17'd54746: data = 8'he9;
      17'd54747: data = 8'hec;
      17'd54748: data = 8'hf1;
      17'd54749: data = 8'hf9;
      17'd54750: data = 8'h01;
      17'd54751: data = 8'h04;
      17'd54752: data = 8'h02;
      17'd54753: data = 8'hfc;
      17'd54754: data = 8'hf2;
      17'd54755: data = 8'hef;
      17'd54756: data = 8'he9;
      17'd54757: data = 8'he7;
      17'd54758: data = 8'he7;
      17'd54759: data = 8'hef;
      17'd54760: data = 8'hef;
      17'd54761: data = 8'he7;
      17'd54762: data = 8'he3;
      17'd54763: data = 8'he4;
      17'd54764: data = 8'hd8;
      17'd54765: data = 8'hd1;
      17'd54766: data = 8'hd5;
      17'd54767: data = 8'hd5;
      17'd54768: data = 8'heb;
      17'd54769: data = 8'hfa;
      17'd54770: data = 8'hfc;
      17'd54771: data = 8'h00;
      17'd54772: data = 8'hf9;
      17'd54773: data = 8'he2;
      17'd54774: data = 8'hcd;
      17'd54775: data = 8'hc1;
      17'd54776: data = 8'hc0;
      17'd54777: data = 8'hce;
      17'd54778: data = 8'he7;
      17'd54779: data = 8'hf5;
      17'd54780: data = 8'h00;
      17'd54781: data = 8'hf9;
      17'd54782: data = 8'hec;
      17'd54783: data = 8'he5;
      17'd54784: data = 8'he5;
      17'd54785: data = 8'hf4;
      17'd54786: data = 8'hfa;
      17'd54787: data = 8'hfd;
      17'd54788: data = 8'hfc;
      17'd54789: data = 8'he7;
      17'd54790: data = 8'hd5;
      17'd54791: data = 8'hcb;
      17'd54792: data = 8'hcb;
      17'd54793: data = 8'hde;
      17'd54794: data = 8'hef;
      17'd54795: data = 8'hf6;
      17'd54796: data = 8'hfa;
      17'd54797: data = 8'hf5;
      17'd54798: data = 8'hec;
      17'd54799: data = 8'he7;
      17'd54800: data = 8'he7;
      17'd54801: data = 8'hed;
      17'd54802: data = 8'hfc;
      17'd54803: data = 8'hfa;
      17'd54804: data = 8'hf5;
      17'd54805: data = 8'hf1;
      17'd54806: data = 8'he5;
      17'd54807: data = 8'he7;
      17'd54808: data = 8'he7;
      17'd54809: data = 8'hf6;
      17'd54810: data = 8'h0c;
      17'd54811: data = 8'h16;
      17'd54812: data = 8'h1c;
      17'd54813: data = 8'h1b;
      17'd54814: data = 8'h12;
      17'd54815: data = 8'h0c;
      17'd54816: data = 8'h0c;
      17'd54817: data = 8'h0e;
      17'd54818: data = 8'h19;
      17'd54819: data = 8'h1b;
      17'd54820: data = 8'h1b;
      17'd54821: data = 8'h1c;
      17'd54822: data = 8'h1a;
      17'd54823: data = 8'h13;
      17'd54824: data = 8'h1f;
      17'd54825: data = 8'h26;
      17'd54826: data = 8'h2d;
      17'd54827: data = 8'h3a;
      17'd54828: data = 8'h39;
      17'd54829: data = 8'h31;
      17'd54830: data = 8'h1c;
      17'd54831: data = 8'h1c;
      17'd54832: data = 8'h1a;
      17'd54833: data = 8'h23;
      17'd54834: data = 8'h24;
      17'd54835: data = 8'h26;
      17'd54836: data = 8'h22;
      17'd54837: data = 8'h11;
      17'd54838: data = 8'h09;
      17'd54839: data = 8'h05;
      17'd54840: data = 8'h11;
      17'd54841: data = 8'h19;
      17'd54842: data = 8'h27;
      17'd54843: data = 8'h24;
      17'd54844: data = 8'h19;
      17'd54845: data = 8'h00;
      17'd54846: data = 8'hfc;
      17'd54847: data = 8'hf1;
      17'd54848: data = 8'hec;
      17'd54849: data = 8'h02;
      17'd54850: data = 8'h09;
      17'd54851: data = 8'h01;
      17'd54852: data = 8'hf5;
      17'd54853: data = 8'he9;
      17'd54854: data = 8'he7;
      17'd54855: data = 8'he5;
      17'd54856: data = 8'h01;
      17'd54857: data = 8'h0c;
      17'd54858: data = 8'h13;
      17'd54859: data = 8'h0a;
      17'd54860: data = 8'he0;
      17'd54861: data = 8'hd5;
      17'd54862: data = 8'hb5;
      17'd54863: data = 8'hb3;
      17'd54864: data = 8'hc1;
      17'd54865: data = 8'hd3;
      17'd54866: data = 8'hec;
      17'd54867: data = 8'he9;
      17'd54868: data = 8'hec;
      17'd54869: data = 8'he4;
      17'd54870: data = 8'hed;
      17'd54871: data = 8'h01;
      17'd54872: data = 8'h1f;
      17'd54873: data = 8'h43;
      17'd54874: data = 8'h40;
      17'd54875: data = 8'h3c;
      17'd54876: data = 8'h2c;
      17'd54877: data = 8'h0d;
      17'd54878: data = 8'h06;
      17'd54879: data = 8'h0e;
      17'd54880: data = 8'h1b;
      17'd54881: data = 8'h2b;
      17'd54882: data = 8'h23;
      17'd54883: data = 8'h23;
      17'd54884: data = 8'h1f;
      17'd54885: data = 8'h23;
      17'd54886: data = 8'h39;
      17'd54887: data = 8'h5a;
      17'd54888: data = 8'h6a;
      17'd54889: data = 8'h68;
      17'd54890: data = 8'h5a;
      17'd54891: data = 8'h3c;
      17'd54892: data = 8'h23;
      17'd54893: data = 8'h1c;
      17'd54894: data = 8'h1c;
      17'd54895: data = 8'h29;
      17'd54896: data = 8'h24;
      17'd54897: data = 8'h0d;
      17'd54898: data = 8'h00;
      17'd54899: data = 8'he5;
      17'd54900: data = 8'he0;
      17'd54901: data = 8'hf1;
      17'd54902: data = 8'h05;
      17'd54903: data = 8'h13;
      17'd54904: data = 8'h0c;
      17'd54905: data = 8'hfd;
      17'd54906: data = 8'he4;
      17'd54907: data = 8'hcd;
      17'd54908: data = 8'hc4;
      17'd54909: data = 8'hc1;
      17'd54910: data = 8'hc6;
      17'd54911: data = 8'hb4;
      17'd54912: data = 8'ha4;
      17'd54913: data = 8'h97;
      17'd54914: data = 8'h8c;
      17'd54915: data = 8'h97;
      17'd54916: data = 8'ha8;
      17'd54917: data = 8'hc4;
      17'd54918: data = 8'hd3;
      17'd54919: data = 8'hce;
      17'd54920: data = 8'hcb;
      17'd54921: data = 8'hc9;
      17'd54922: data = 8'hcb;
      17'd54923: data = 8'hd2;
      17'd54924: data = 8'he4;
      17'd54925: data = 8'hec;
      17'd54926: data = 8'he3;
      17'd54927: data = 8'hdb;
      17'd54928: data = 8'hd3;
      17'd54929: data = 8'hda;
      17'd54930: data = 8'heb;
      17'd54931: data = 8'h04;
      17'd54932: data = 8'h26;
      17'd54933: data = 8'h35;
      17'd54934: data = 8'h3c;
      17'd54935: data = 8'h46;
      17'd54936: data = 8'h4e;
      17'd54937: data = 8'h5a;
      17'd54938: data = 8'h63;
      17'd54939: data = 8'h6a;
      17'd54940: data = 8'h60;
      17'd54941: data = 8'h52;
      17'd54942: data = 8'h46;
      17'd54943: data = 8'h3c;
      17'd54944: data = 8'h42;
      17'd54945: data = 8'h4a;
      17'd54946: data = 8'h52;
      17'd54947: data = 8'h57;
      17'd54948: data = 8'h4d;
      17'd54949: data = 8'h46;
      17'd54950: data = 8'h43;
      17'd54951: data = 8'h45;
      17'd54952: data = 8'h4d;
      17'd54953: data = 8'h4d;
      17'd54954: data = 8'h47;
      17'd54955: data = 8'h34;
      17'd54956: data = 8'h13;
      17'd54957: data = 8'hf9;
      17'd54958: data = 8'he7;
      17'd54959: data = 8'hde;
      17'd54960: data = 8'hda;
      17'd54961: data = 8'hd8;
      17'd54962: data = 8'hd1;
      17'd54963: data = 8'hc5;
      17'd54964: data = 8'hbd;
      17'd54965: data = 8'hb8;
      17'd54966: data = 8'hb9;
      17'd54967: data = 8'hbd;
      17'd54968: data = 8'hc2;
      17'd54969: data = 8'hc2;
      17'd54970: data = 8'hb4;
      17'd54971: data = 8'ha6;
      17'd54972: data = 8'h9f;
      17'd54973: data = 8'h97;
      17'd54974: data = 8'h97;
      17'd54975: data = 8'h9b;
      17'd54976: data = 8'ha3;
      17'd54977: data = 8'haa;
      17'd54978: data = 8'hb0;
      17'd54979: data = 8'hbc;
      17'd54980: data = 8'hcb;
      17'd54981: data = 8'he0;
      17'd54982: data = 8'he4;
      17'd54983: data = 8'hec;
      17'd54984: data = 8'hf5;
      17'd54985: data = 8'hf5;
      17'd54986: data = 8'hfc;
      17'd54987: data = 8'h09;
      17'd54988: data = 8'h11;
      17'd54989: data = 8'h12;
      17'd54990: data = 8'h15;
      17'd54991: data = 8'h15;
      17'd54992: data = 8'h15;
      17'd54993: data = 8'h1e;
      17'd54994: data = 8'h27;
      17'd54995: data = 8'h34;
      17'd54996: data = 8'h39;
      17'd54997: data = 8'h3c;
      17'd54998: data = 8'h40;
      17'd54999: data = 8'h3d;
      17'd55000: data = 8'h3d;
      17'd55001: data = 8'h39;
      17'd55002: data = 8'h33;
      17'd55003: data = 8'h2b;
      17'd55004: data = 8'h1e;
      17'd55005: data = 8'h13;
      17'd55006: data = 8'h0e;
      17'd55007: data = 8'h0c;
      17'd55008: data = 8'h09;
      17'd55009: data = 8'h06;
      17'd55010: data = 8'h00;
      17'd55011: data = 8'hf2;
      17'd55012: data = 8'he7;
      17'd55013: data = 8'hdc;
      17'd55014: data = 8'hd8;
      17'd55015: data = 8'hd8;
      17'd55016: data = 8'hd6;
      17'd55017: data = 8'hd1;
      17'd55018: data = 8'hc4;
      17'd55019: data = 8'hb8;
      17'd55020: data = 8'hac;
      17'd55021: data = 8'ha8;
      17'd55022: data = 8'ha8;
      17'd55023: data = 8'hae;
      17'd55024: data = 8'hb3;
      17'd55025: data = 8'hb3;
      17'd55026: data = 8'hb5;
      17'd55027: data = 8'hb5;
      17'd55028: data = 8'hb3;
      17'd55029: data = 8'hb8;
      17'd55030: data = 8'hbb;
      17'd55031: data = 8'hc0;
      17'd55032: data = 8'hc6;
      17'd55033: data = 8'hcd;
      17'd55034: data = 8'hd1;
      17'd55035: data = 8'hd5;
      17'd55036: data = 8'he0;
      17'd55037: data = 8'heb;
      17'd55038: data = 8'hf5;
      17'd55039: data = 8'h01;
      17'd55040: data = 8'h0c;
      17'd55041: data = 8'h12;
      17'd55042: data = 8'h15;
      17'd55043: data = 8'h1c;
      17'd55044: data = 8'h27;
      17'd55045: data = 8'h31;
      17'd55046: data = 8'h34;
      17'd55047: data = 8'h39;
      17'd55048: data = 8'h33;
      17'd55049: data = 8'h33;
      17'd55050: data = 8'h3e;
      17'd55051: data = 8'h3d;
      17'd55052: data = 8'h4a;
      17'd55053: data = 8'h4b;
      17'd55054: data = 8'h4d;
      17'd55055: data = 8'h4d;
      17'd55056: data = 8'h46;
      17'd55057: data = 8'h3e;
      17'd55058: data = 8'h39;
      17'd55059: data = 8'h24;
      17'd55060: data = 8'h31;
      17'd55061: data = 8'h2f;
      17'd55062: data = 8'h12;
      17'd55063: data = 8'h26;
      17'd55064: data = 8'h12;
      17'd55065: data = 8'h06;
      17'd55066: data = 8'hfd;
      17'd55067: data = 8'hf6;
      17'd55068: data = 8'hf5;
      17'd55069: data = 8'hfc;
      17'd55070: data = 8'he7;
      17'd55071: data = 8'he9;
      17'd55072: data = 8'hf1;
      17'd55073: data = 8'hdc;
      17'd55074: data = 8'hde;
      17'd55075: data = 8'hec;
      17'd55076: data = 8'hd6;
      17'd55077: data = 8'hcb;
      17'd55078: data = 8'hd1;
      17'd55079: data = 8'hc2;
      17'd55080: data = 8'hd3;
      17'd55081: data = 8'hda;
      17'd55082: data = 8'he3;
      17'd55083: data = 8'hf9;
      17'd55084: data = 8'hef;
      17'd55085: data = 8'hd3;
      17'd55086: data = 8'hec;
      17'd55087: data = 8'hed;
      17'd55088: data = 8'heb;
      17'd55089: data = 8'h09;
      17'd55090: data = 8'h0c;
      17'd55091: data = 8'h26;
      17'd55092: data = 8'h2f;
      17'd55093: data = 8'h24;
      17'd55094: data = 8'h1e;
      17'd55095: data = 8'h05;
      17'd55096: data = 8'hde;
      17'd55097: data = 8'he2;
      17'd55098: data = 8'he5;
      17'd55099: data = 8'he0;
      17'd55100: data = 8'h09;
      17'd55101: data = 8'h1e;
      17'd55102: data = 8'h26;
      17'd55103: data = 8'h40;
      17'd55104: data = 8'h3e;
      17'd55105: data = 8'h46;
      17'd55106: data = 8'h54;
      17'd55107: data = 8'h4a;
      17'd55108: data = 8'h5c;
      17'd55109: data = 8'h5d;
      17'd55110: data = 8'h3e;
      17'd55111: data = 8'h39;
      17'd55112: data = 8'h2d;
      17'd55113: data = 8'h1e;
      17'd55114: data = 8'h11;
      17'd55115: data = 8'h19;
      17'd55116: data = 8'h06;
      17'd55117: data = 8'h0d;
      17'd55118: data = 8'h0e;
      17'd55119: data = 8'h15;
      17'd55120: data = 8'h43;
      17'd55121: data = 8'h40;
      17'd55122: data = 8'h4a;
      17'd55123: data = 8'h4e;
      17'd55124: data = 8'h29;
      17'd55125: data = 8'h01;
      17'd55126: data = 8'hec;
      17'd55127: data = 8'hd3;
      17'd55128: data = 8'hd1;
      17'd55129: data = 8'hd2;
      17'd55130: data = 8'hd2;
      17'd55131: data = 8'hd2;
      17'd55132: data = 8'hca;
      17'd55133: data = 8'hbc;
      17'd55134: data = 8'hc5;
      17'd55135: data = 8'hd3;
      17'd55136: data = 8'hd3;
      17'd55137: data = 8'he7;
      17'd55138: data = 8'he5;
      17'd55139: data = 8'hdb;
      17'd55140: data = 8'hdc;
      17'd55141: data = 8'hcd;
      17'd55142: data = 8'hc5;
      17'd55143: data = 8'hbb;
      17'd55144: data = 8'ha8;
      17'd55145: data = 8'h9d;
      17'd55146: data = 8'h9b;
      17'd55147: data = 8'ha1;
      17'd55148: data = 8'hae;
      17'd55149: data = 8'hcd;
      17'd55150: data = 8'he5;
      17'd55151: data = 8'h00;
      17'd55152: data = 8'h15;
      17'd55153: data = 8'h19;
      17'd55154: data = 8'h1a;
      17'd55155: data = 8'h13;
      17'd55156: data = 8'h0e;
      17'd55157: data = 8'h11;
      17'd55158: data = 8'h0d;
      17'd55159: data = 8'h0d;
      17'd55160: data = 8'h11;
      17'd55161: data = 8'h16;
      17'd55162: data = 8'h16;
      17'd55163: data = 8'h22;
      17'd55164: data = 8'h2f;
      17'd55165: data = 8'h36;
      17'd55166: data = 8'h4d;
      17'd55167: data = 8'h5d;
      17'd55168: data = 8'h6a;
      17'd55169: data = 8'h74;
      17'd55170: data = 8'h70;
      17'd55171: data = 8'h68;
      17'd55172: data = 8'h5c;
      17'd55173: data = 8'h46;
      17'd55174: data = 8'h36;
      17'd55175: data = 8'h29;
      17'd55176: data = 8'h1b;
      17'd55177: data = 8'h16;
      17'd55178: data = 8'h1a;
      17'd55179: data = 8'h1f;
      17'd55180: data = 8'h29;
      17'd55181: data = 8'h2d;
      17'd55182: data = 8'h2c;
      17'd55183: data = 8'h2b;
      17'd55184: data = 8'h1c;
      17'd55185: data = 8'h12;
      17'd55186: data = 8'h05;
      17'd55187: data = 8'hf6;
      17'd55188: data = 8'hec;
      17'd55189: data = 8'he0;
      17'd55190: data = 8'hd3;
      17'd55191: data = 8'hc1;
      17'd55192: data = 8'hb5;
      17'd55193: data = 8'hab;
      17'd55194: data = 8'haa;
      17'd55195: data = 8'hb1;
      17'd55196: data = 8'hbb;
      17'd55197: data = 8'hca;
      17'd55198: data = 8'hd5;
      17'd55199: data = 8'hda;
      17'd55200: data = 8'hd8;
      17'd55201: data = 8'hd6;
      17'd55202: data = 8'hce;
      17'd55203: data = 8'hc9;
      17'd55204: data = 8'hc1;
      17'd55205: data = 8'hbc;
      17'd55206: data = 8'hbb;
      17'd55207: data = 8'hbb;
      17'd55208: data = 8'hc6;
      17'd55209: data = 8'hd3;
      17'd55210: data = 8'he3;
      17'd55211: data = 8'hf1;
      17'd55212: data = 8'hfd;
      17'd55213: data = 8'h05;
      17'd55214: data = 8'h0e;
      17'd55215: data = 8'h1a;
      17'd55216: data = 8'h24;
      17'd55217: data = 8'h26;
      17'd55218: data = 8'h23;
      17'd55219: data = 8'h22;
      17'd55220: data = 8'h1b;
      17'd55221: data = 8'h15;
      17'd55222: data = 8'h0e;
      17'd55223: data = 8'h11;
      17'd55224: data = 8'h12;
      17'd55225: data = 8'h16;
      17'd55226: data = 8'h22;
      17'd55227: data = 8'h27;
      17'd55228: data = 8'h2c;
      17'd55229: data = 8'h2b;
      17'd55230: data = 8'h27;
      17'd55231: data = 8'h1e;
      17'd55232: data = 8'h11;
      17'd55233: data = 8'h04;
      17'd55234: data = 8'hf6;
      17'd55235: data = 8'hf1;
      17'd55236: data = 8'he5;
      17'd55237: data = 8'hde;
      17'd55238: data = 8'hde;
      17'd55239: data = 8'hda;
      17'd55240: data = 8'hd5;
      17'd55241: data = 8'hd5;
      17'd55242: data = 8'hd3;
      17'd55243: data = 8'hd1;
      17'd55244: data = 8'hd2;
      17'd55245: data = 8'hd2;
      17'd55246: data = 8'hce;
      17'd55247: data = 8'hca;
      17'd55248: data = 8'hc4;
      17'd55249: data = 8'hbd;
      17'd55250: data = 8'hb9;
      17'd55251: data = 8'hb3;
      17'd55252: data = 8'hb1;
      17'd55253: data = 8'hb9;
      17'd55254: data = 8'hbc;
      17'd55255: data = 8'hc4;
      17'd55256: data = 8'hd3;
      17'd55257: data = 8'he2;
      17'd55258: data = 8'he4;
      17'd55259: data = 8'heb;
      17'd55260: data = 8'hf1;
      17'd55261: data = 8'hec;
      17'd55262: data = 8'hec;
      17'd55263: data = 8'heb;
      17'd55264: data = 8'hf2;
      17'd55265: data = 8'hf5;
      17'd55266: data = 8'hfa;
      17'd55267: data = 8'h06;
      17'd55268: data = 8'h0a;
      17'd55269: data = 8'h0c;
      17'd55270: data = 8'h15;
      17'd55271: data = 8'h1a;
      17'd55272: data = 8'h1c;
      17'd55273: data = 8'h2c;
      17'd55274: data = 8'h2b;
      17'd55275: data = 8'h2c;
      17'd55276: data = 8'h34;
      17'd55277: data = 8'h2d;
      17'd55278: data = 8'h29;
      17'd55279: data = 8'h24;
      17'd55280: data = 8'h1f;
      17'd55281: data = 8'h2d;
      17'd55282: data = 8'h1f;
      17'd55283: data = 8'h19;
      17'd55284: data = 8'h27;
      17'd55285: data = 8'h15;
      17'd55286: data = 8'h13;
      17'd55287: data = 8'h1f;
      17'd55288: data = 8'h1b;
      17'd55289: data = 8'h13;
      17'd55290: data = 8'h05;
      17'd55291: data = 8'h02;
      17'd55292: data = 8'hfd;
      17'd55293: data = 8'hfc;
      17'd55294: data = 8'hf9;
      17'd55295: data = 8'hfe;
      17'd55296: data = 8'hed;
      17'd55297: data = 8'hef;
      17'd55298: data = 8'hec;
      17'd55299: data = 8'hd8;
      17'd55300: data = 8'hfe;
      17'd55301: data = 8'he9;
      17'd55302: data = 8'hf4;
      17'd55303: data = 8'hfa;
      17'd55304: data = 8'hf2;
      17'd55305: data = 8'hec;
      17'd55306: data = 8'he5;
      17'd55307: data = 8'hfd;
      17'd55308: data = 8'he3;
      17'd55309: data = 8'hf9;
      17'd55310: data = 8'hf6;
      17'd55311: data = 8'hf9;
      17'd55312: data = 8'h00;
      17'd55313: data = 8'hf5;
      17'd55314: data = 8'h1b;
      17'd55315: data = 8'h12;
      17'd55316: data = 8'h1b;
      17'd55317: data = 8'h1f;
      17'd55318: data = 8'h1f;
      17'd55319: data = 8'h27;
      17'd55320: data = 8'h22;
      17'd55321: data = 8'h39;
      17'd55322: data = 8'h31;
      17'd55323: data = 8'h2f;
      17'd55324: data = 8'h2d;
      17'd55325: data = 8'h09;
      17'd55326: data = 8'hf4;
      17'd55327: data = 8'hfc;
      17'd55328: data = 8'h05;
      17'd55329: data = 8'hef;
      17'd55330: data = 8'hf2;
      17'd55331: data = 8'h09;
      17'd55332: data = 8'h01;
      17'd55333: data = 8'h02;
      17'd55334: data = 8'h1e;
      17'd55335: data = 8'h4b;
      17'd55336: data = 8'h5b;
      17'd55337: data = 8'h45;
      17'd55338: data = 8'h40;
      17'd55339: data = 8'h2c;
      17'd55340: data = 8'hfc;
      17'd55341: data = 8'hf1;
      17'd55342: data = 8'hfd;
      17'd55343: data = 8'h0d;
      17'd55344: data = 8'h06;
      17'd55345: data = 8'h00;
      17'd55346: data = 8'hfa;
      17'd55347: data = 8'hef;
      17'd55348: data = 8'h01;
      17'd55349: data = 8'h0e;
      17'd55350: data = 8'h29;
      17'd55351: data = 8'h2d;
      17'd55352: data = 8'h2d;
      17'd55353: data = 8'h27;
      17'd55354: data = 8'h02;
      17'd55355: data = 8'h06;
      17'd55356: data = 8'h04;
      17'd55357: data = 8'hfe;
      17'd55358: data = 8'hef;
      17'd55359: data = 8'hd8;
      17'd55360: data = 8'hd1;
      17'd55361: data = 8'hb9;
      17'd55362: data = 8'hbc;
      17'd55363: data = 8'hda;
      17'd55364: data = 8'h0c;
      17'd55365: data = 8'h16;
      17'd55366: data = 8'h12;
      17'd55367: data = 8'h1c;
      17'd55368: data = 8'h00;
      17'd55369: data = 8'he5;
      17'd55370: data = 8'hdb;
      17'd55371: data = 8'he2;
      17'd55372: data = 8'heb;
      17'd55373: data = 8'hd3;
      17'd55374: data = 8'hd1;
      17'd55375: data = 8'hd6;
      17'd55376: data = 8'hc4;
      17'd55377: data = 8'hc6;
      17'd55378: data = 8'hd3;
      17'd55379: data = 8'he5;
      17'd55380: data = 8'hf2;
      17'd55381: data = 8'h01;
      17'd55382: data = 8'h05;
      17'd55383: data = 8'h0a;
      17'd55384: data = 8'h16;
      17'd55385: data = 8'h11;
      17'd55386: data = 8'h19;
      17'd55387: data = 8'h0e;
      17'd55388: data = 8'hfd;
      17'd55389: data = 8'hfa;
      17'd55390: data = 8'he9;
      17'd55391: data = 8'hec;
      17'd55392: data = 8'hfd;
      17'd55393: data = 8'h0e;
      17'd55394: data = 8'h22;
      17'd55395: data = 8'h35;
      17'd55396: data = 8'h46;
      17'd55397: data = 8'h4a;
      17'd55398: data = 8'h4a;
      17'd55399: data = 8'h3a;
      17'd55400: data = 8'h40;
      17'd55401: data = 8'h39;
      17'd55402: data = 8'h29;
      17'd55403: data = 8'h2b;
      17'd55404: data = 8'h29;
      17'd55405: data = 8'h1f;
      17'd55406: data = 8'h12;
      17'd55407: data = 8'h11;
      17'd55408: data = 8'h12;
      17'd55409: data = 8'h16;
      17'd55410: data = 8'h1c;
      17'd55411: data = 8'h26;
      17'd55412: data = 8'h2d;
      17'd55413: data = 8'h27;
      17'd55414: data = 8'h24;
      17'd55415: data = 8'h1f;
      17'd55416: data = 8'h19;
      17'd55417: data = 8'h0e;
      17'd55418: data = 8'hfc;
      17'd55419: data = 8'he9;
      17'd55420: data = 8'hda;
      17'd55421: data = 8'hcb;
      17'd55422: data = 8'hc6;
      17'd55423: data = 8'hcd;
      17'd55424: data = 8'hdc;
      17'd55425: data = 8'he7;
      17'd55426: data = 8'he7;
      17'd55427: data = 8'he7;
      17'd55428: data = 8'he0;
      17'd55429: data = 8'he4;
      17'd55430: data = 8'he4;
      17'd55431: data = 8'he4;
      17'd55432: data = 8'he7;
      17'd55433: data = 8'he3;
      17'd55434: data = 8'hdb;
      17'd55435: data = 8'hce;
      17'd55436: data = 8'hce;
      17'd55437: data = 8'hd1;
      17'd55438: data = 8'hd3;
      17'd55439: data = 8'hdb;
      17'd55440: data = 8'he7;
      17'd55441: data = 8'hf5;
      17'd55442: data = 8'hf6;
      17'd55443: data = 8'hfd;
      17'd55444: data = 8'h06;
      17'd55445: data = 8'h0e;
      17'd55446: data = 8'h0e;
      17'd55447: data = 8'h0e;
      17'd55448: data = 8'h0a;
      17'd55449: data = 8'h01;
      17'd55450: data = 8'hfa;
      17'd55451: data = 8'hf6;
      17'd55452: data = 8'hfc;
      17'd55453: data = 8'h02;
      17'd55454: data = 8'h06;
      17'd55455: data = 8'h09;
      17'd55456: data = 8'h0a;
      17'd55457: data = 8'h0c;
      17'd55458: data = 8'h0e;
      17'd55459: data = 8'h11;
      17'd55460: data = 8'h11;
      17'd55461: data = 8'h0e;
      17'd55462: data = 8'h06;
      17'd55463: data = 8'hfd;
      17'd55464: data = 8'hf1;
      17'd55465: data = 8'he9;
      17'd55466: data = 8'he5;
      17'd55467: data = 8'he3;
      17'd55468: data = 8'hdc;
      17'd55469: data = 8'hda;
      17'd55470: data = 8'hdb;
      17'd55471: data = 8'hd5;
      17'd55472: data = 8'hdb;
      17'd55473: data = 8'he0;
      17'd55474: data = 8'hde;
      17'd55475: data = 8'hdb;
      17'd55476: data = 8'hd8;
      17'd55477: data = 8'hd5;
      17'd55478: data = 8'hcd;
      17'd55479: data = 8'hca;
      17'd55480: data = 8'hc5;
      17'd55481: data = 8'hcb;
      17'd55482: data = 8'hcb;
      17'd55483: data = 8'hc9;
      17'd55484: data = 8'hd2;
      17'd55485: data = 8'hd8;
      17'd55486: data = 8'he0;
      17'd55487: data = 8'he9;
      17'd55488: data = 8'hf1;
      17'd55489: data = 8'hf4;
      17'd55490: data = 8'hf1;
      17'd55491: data = 8'hed;
      17'd55492: data = 8'hed;
      17'd55493: data = 8'hf1;
      17'd55494: data = 8'hf4;
      17'd55495: data = 8'hf9;
      17'd55496: data = 8'hfa;
      17'd55497: data = 8'hfa;
      17'd55498: data = 8'hf9;
      17'd55499: data = 8'hfa;
      17'd55500: data = 8'hfe;
      17'd55501: data = 8'h0e;
      17'd55502: data = 8'h1e;
      17'd55503: data = 8'h1e;
      17'd55504: data = 8'h1e;
      17'd55505: data = 8'h1a;
      17'd55506: data = 8'h11;
      17'd55507: data = 8'h13;
      17'd55508: data = 8'h15;
      17'd55509: data = 8'h12;
      17'd55510: data = 8'h1f;
      17'd55511: data = 8'h12;
      17'd55512: data = 8'h0e;
      17'd55513: data = 8'h15;
      17'd55514: data = 8'h05;
      17'd55515: data = 8'h16;
      17'd55516: data = 8'h1b;
      17'd55517: data = 8'h06;
      17'd55518: data = 8'h1b;
      17'd55519: data = 8'h15;
      17'd55520: data = 8'hf5;
      17'd55521: data = 8'h04;
      17'd55522: data = 8'h0a;
      17'd55523: data = 8'h00;
      17'd55524: data = 8'hfc;
      17'd55525: data = 8'heb;
      17'd55526: data = 8'hf2;
      17'd55527: data = 8'he7;
      17'd55528: data = 8'hef;
      17'd55529: data = 8'hfd;
      17'd55530: data = 8'hf1;
      17'd55531: data = 8'hf1;
      17'd55532: data = 8'hfa;
      17'd55533: data = 8'hf5;
      17'd55534: data = 8'hf6;
      17'd55535: data = 8'h00;
      17'd55536: data = 8'hf1;
      17'd55537: data = 8'h05;
      17'd55538: data = 8'hf9;
      17'd55539: data = 8'hfc;
      17'd55540: data = 8'h04;
      17'd55541: data = 8'hf1;
      17'd55542: data = 8'h09;
      17'd55543: data = 8'h0c;
      17'd55544: data = 8'h02;
      17'd55545: data = 8'h1b;
      17'd55546: data = 8'h11;
      17'd55547: data = 8'h04;
      17'd55548: data = 8'h19;
      17'd55549: data = 8'h1f;
      17'd55550: data = 8'h2d;
      17'd55551: data = 8'h4f;
      17'd55552: data = 8'h3e;
      17'd55553: data = 8'h24;
      17'd55554: data = 8'h1b;
      17'd55555: data = 8'heb;
      17'd55556: data = 8'hb3;
      17'd55557: data = 8'hc5;
      17'd55558: data = 8'he3;
      17'd55559: data = 8'hf2;
      17'd55560: data = 8'h13;
      17'd55561: data = 8'h31;
      17'd55562: data = 8'h45;
      17'd55563: data = 8'h42;
      17'd55564: data = 8'h3d;
      17'd55565: data = 8'h5a;
      17'd55566: data = 8'h4a;
      17'd55567: data = 8'h2b;
      17'd55568: data = 8'h26;
      17'd55569: data = 8'h06;
      17'd55570: data = 8'hde;
      17'd55571: data = 8'hf6;
      17'd55572: data = 8'h09;
      17'd55573: data = 8'hf9;
      17'd55574: data = 8'h1a;
      17'd55575: data = 8'h19;
      17'd55576: data = 8'h02;
      17'd55577: data = 8'hfe;
      17'd55578: data = 8'hfd;
      17'd55579: data = 8'h1b;
      17'd55580: data = 8'h39;
      17'd55581: data = 8'h40;
      17'd55582: data = 8'h4e;
      17'd55583: data = 8'h35;
      17'd55584: data = 8'hfd;
      17'd55585: data = 8'he0;
      17'd55586: data = 8'hc2;
      17'd55587: data = 8'hbd;
      17'd55588: data = 8'hcd;
      17'd55589: data = 8'hc4;
      17'd55590: data = 8'hd2;
      17'd55591: data = 8'he9;
      17'd55592: data = 8'he3;
      17'd55593: data = 8'hed;
      17'd55594: data = 8'h15;
      17'd55595: data = 8'h11;
      17'd55596: data = 8'h00;
      17'd55597: data = 8'hf9;
      17'd55598: data = 8'hd6;
      17'd55599: data = 8'hc4;
      17'd55600: data = 8'hbb;
      17'd55601: data = 8'hc5;
      17'd55602: data = 8'hd8;
      17'd55603: data = 8'hd5;
      17'd55604: data = 8'hd6;
      17'd55605: data = 8'hd5;
      17'd55606: data = 8'hbc;
      17'd55607: data = 8'hc5;
      17'd55608: data = 8'he7;
      17'd55609: data = 8'hfa;
      17'd55610: data = 8'h15;
      17'd55611: data = 8'h31;
      17'd55612: data = 8'h29;
      17'd55613: data = 8'h1f;
      17'd55614: data = 8'h1a;
      17'd55615: data = 8'h09;
      17'd55616: data = 8'h0a;
      17'd55617: data = 8'h01;
      17'd55618: data = 8'hf4;
      17'd55619: data = 8'h02;
      17'd55620: data = 8'h05;
      17'd55621: data = 8'h12;
      17'd55622: data = 8'h2d;
      17'd55623: data = 8'h42;
      17'd55624: data = 8'h5a;
      17'd55625: data = 8'h5c;
      17'd55626: data = 8'h4f;
      17'd55627: data = 8'h4a;
      17'd55628: data = 8'h3c;
      17'd55629: data = 8'h27;
      17'd55630: data = 8'h33;
      17'd55631: data = 8'h34;
      17'd55632: data = 8'h27;
      17'd55633: data = 8'h2c;
      17'd55634: data = 8'h1e;
      17'd55635: data = 8'h0a;
      17'd55636: data = 8'h0a;
      17'd55637: data = 8'h06;
      17'd55638: data = 8'h0a;
      17'd55639: data = 8'h16;
      17'd55640: data = 8'h1c;
      17'd55641: data = 8'h24;
      17'd55642: data = 8'h24;
      17'd55643: data = 8'h19;
      17'd55644: data = 8'h13;
      17'd55645: data = 8'h00;
      17'd55646: data = 8'heb;
      17'd55647: data = 8'hde;
      17'd55648: data = 8'hce;
      17'd55649: data = 8'hc0;
      17'd55650: data = 8'hbd;
      17'd55651: data = 8'hc2;
      17'd55652: data = 8'hd1;
      17'd55653: data = 8'he5;
      17'd55654: data = 8'he7;
      17'd55655: data = 8'hec;
      17'd55656: data = 8'hef;
      17'd55657: data = 8'he3;
      17'd55658: data = 8'hde;
      17'd55659: data = 8'he4;
      17'd55660: data = 8'he7;
      17'd55661: data = 8'he9;
      17'd55662: data = 8'he9;
      17'd55663: data = 8'he4;
      17'd55664: data = 8'hdb;
      17'd55665: data = 8'hd6;
      17'd55666: data = 8'hdb;
      17'd55667: data = 8'he7;
      17'd55668: data = 8'hf1;
      17'd55669: data = 8'h01;
      17'd55670: data = 8'h12;
      17'd55671: data = 8'h12;
      17'd55672: data = 8'h1f;
      17'd55673: data = 8'h2c;
      17'd55674: data = 8'h26;
      17'd55675: data = 8'h23;
      17'd55676: data = 8'h1c;
      17'd55677: data = 8'h0a;
      17'd55678: data = 8'hfd;
      17'd55679: data = 8'hf6;
      17'd55680: data = 8'hfc;
      17'd55681: data = 8'h06;
      17'd55682: data = 8'h11;
      17'd55683: data = 8'h19;
      17'd55684: data = 8'h1b;
      17'd55685: data = 8'h1a;
      17'd55686: data = 8'h11;
      17'd55687: data = 8'h0e;
      17'd55688: data = 8'h09;
      17'd55689: data = 8'h02;
      17'd55690: data = 8'hf9;
      17'd55691: data = 8'hed;
      17'd55692: data = 8'he5;
      17'd55693: data = 8'hdb;
      17'd55694: data = 8'hd3;
      17'd55695: data = 8'hd1;
      17'd55696: data = 8'hcd;
      17'd55697: data = 8'hc6;
      17'd55698: data = 8'hca;
      17'd55699: data = 8'hca;
      17'd55700: data = 8'hce;
      17'd55701: data = 8'hd8;
      17'd55702: data = 8'hdc;
      17'd55703: data = 8'hdc;
      17'd55704: data = 8'hd8;
      17'd55705: data = 8'hd1;
      17'd55706: data = 8'hc2;
      17'd55707: data = 8'hb9;
      17'd55708: data = 8'hb8;
      17'd55709: data = 8'hbd;
      17'd55710: data = 8'hc4;
      17'd55711: data = 8'hca;
      17'd55712: data = 8'hda;
      17'd55713: data = 8'he2;
      17'd55714: data = 8'he5;
      17'd55715: data = 8'hf1;
      17'd55716: data = 8'hfa;
      17'd55717: data = 8'h00;
      17'd55718: data = 8'hfe;
      17'd55719: data = 8'hfd;
      17'd55720: data = 8'hfc;
      17'd55721: data = 8'hf6;
      17'd55722: data = 8'hf2;
      17'd55723: data = 8'hf9;
      17'd55724: data = 8'h02;
      17'd55725: data = 8'h02;
      17'd55726: data = 8'h04;
      17'd55727: data = 8'h0d;
      17'd55728: data = 8'h11;
      17'd55729: data = 8'h19;
      17'd55730: data = 8'h1b;
      17'd55731: data = 8'h24;
      17'd55732: data = 8'h2b;
      17'd55733: data = 8'h23;
      17'd55734: data = 8'h22;
      17'd55735: data = 8'h1e;
      17'd55736: data = 8'h13;
      17'd55737: data = 8'h09;
      17'd55738: data = 8'h0c;
      17'd55739: data = 8'h06;
      17'd55740: data = 8'h0a;
      17'd55741: data = 8'h09;
      17'd55742: data = 8'h09;
      17'd55743: data = 8'h0a;
      17'd55744: data = 8'h0d;
      17'd55745: data = 8'h0e;
      17'd55746: data = 8'h0e;
      17'd55747: data = 8'h0c;
      17'd55748: data = 8'h02;
      17'd55749: data = 8'hf9;
      17'd55750: data = 8'hf9;
      17'd55751: data = 8'hec;
      17'd55752: data = 8'he2;
      17'd55753: data = 8'hfd;
      17'd55754: data = 8'hed;
      17'd55755: data = 8'he7;
      17'd55756: data = 8'hfa;
      17'd55757: data = 8'hec;
      17'd55758: data = 8'he7;
      17'd55759: data = 8'he9;
      17'd55760: data = 8'hf9;
      17'd55761: data = 8'hf5;
      17'd55762: data = 8'hf1;
      17'd55763: data = 8'hf4;
      17'd55764: data = 8'h06;
      17'd55765: data = 8'he9;
      17'd55766: data = 8'hf1;
      17'd55767: data = 8'h01;
      17'd55768: data = 8'he3;
      17'd55769: data = 8'hfa;
      17'd55770: data = 8'h06;
      17'd55771: data = 8'h05;
      17'd55772: data = 8'h13;
      17'd55773: data = 8'h3a;
      17'd55774: data = 8'h42;
      17'd55775: data = 8'h42;
      17'd55776: data = 8'h3a;
      17'd55777: data = 8'h0e;
      17'd55778: data = 8'hf6;
      17'd55779: data = 8'hc6;
      17'd55780: data = 8'hc1;
      17'd55781: data = 8'hd6;
      17'd55782: data = 8'hf1;
      17'd55783: data = 8'h1a;
      17'd55784: data = 8'h22;
      17'd55785: data = 8'h2d;
      17'd55786: data = 8'h47;
      17'd55787: data = 8'h3d;
      17'd55788: data = 8'h29;
      17'd55789: data = 8'h56;
      17'd55790: data = 8'h5b;
      17'd55791: data = 8'h29;
      17'd55792: data = 8'h27;
      17'd55793: data = 8'h1a;
      17'd55794: data = 8'hfd;
      17'd55795: data = 8'hfd;
      17'd55796: data = 8'h12;
      17'd55797: data = 8'h13;
      17'd55798: data = 8'h15;
      17'd55799: data = 8'h02;
      17'd55800: data = 8'h00;
      17'd55801: data = 8'h05;
      17'd55802: data = 8'h04;
      17'd55803: data = 8'h40;
      17'd55804: data = 8'h42;
      17'd55805: data = 8'h42;
      17'd55806: data = 8'h40;
      17'd55807: data = 8'h11;
      17'd55808: data = 8'he5;
      17'd55809: data = 8'hd1;
      17'd55810: data = 8'hcb;
      17'd55811: data = 8'hca;
      17'd55812: data = 8'hdc;
      17'd55813: data = 8'hd6;
      17'd55814: data = 8'hd8;
      17'd55815: data = 8'he4;
      17'd55816: data = 8'hda;
      17'd55817: data = 8'he4;
      17'd55818: data = 8'hfa;
      17'd55819: data = 8'hfe;
      17'd55820: data = 8'hf1;
      17'd55821: data = 8'hdc;
      17'd55822: data = 8'hd6;
      17'd55823: data = 8'hd6;
      17'd55824: data = 8'hbb;
      17'd55825: data = 8'hd2;
      17'd55826: data = 8'he0;
      17'd55827: data = 8'hc6;
      17'd55828: data = 8'hc5;
      17'd55829: data = 8'hc0;
      17'd55830: data = 8'hc0;
      17'd55831: data = 8'hc5;
      17'd55832: data = 8'heb;
      17'd55833: data = 8'h00;
      17'd55834: data = 8'h19;
      17'd55835: data = 8'h2b;
      17'd55836: data = 8'h1f;
      17'd55837: data = 8'h1c;
      17'd55838: data = 8'h0a;
      17'd55839: data = 8'h09;
      17'd55840: data = 8'h09;
      17'd55841: data = 8'hfe;
      17'd55842: data = 8'h09;
      17'd55843: data = 8'h12;
      17'd55844: data = 8'h16;
      17'd55845: data = 8'h29;
      17'd55846: data = 8'h3a;
      17'd55847: data = 8'h46;
      17'd55848: data = 8'h54;
      17'd55849: data = 8'h4f;
      17'd55850: data = 8'h4d;
      17'd55851: data = 8'h4e;
      17'd55852: data = 8'h46;
      17'd55853: data = 8'h36;
      17'd55854: data = 8'h3d;
      17'd55855: data = 8'h40;
      17'd55856: data = 8'h33;
      17'd55857: data = 8'h31;
      17'd55858: data = 8'h1f;
      17'd55859: data = 8'h1a;
      17'd55860: data = 8'h0c;
      17'd55861: data = 8'h06;
      17'd55862: data = 8'h13;
      17'd55863: data = 8'h19;
      17'd55864: data = 8'h23;
      17'd55865: data = 8'h26;
      17'd55866: data = 8'h1e;
      17'd55867: data = 8'h12;
      17'd55868: data = 8'h06;
      17'd55869: data = 8'hf5;
      17'd55870: data = 8'he3;
      17'd55871: data = 8'he2;
      17'd55872: data = 8'hd5;
      17'd55873: data = 8'hcb;
      17'd55874: data = 8'hc9;
      17'd55875: data = 8'hca;
      17'd55876: data = 8'hd3;
      17'd55877: data = 8'hda;
      17'd55878: data = 8'he0;
      17'd55879: data = 8'he5;
      17'd55880: data = 8'he7;
      17'd55881: data = 8'he5;
      17'd55882: data = 8'he4;
      17'd55883: data = 8'he4;
      17'd55884: data = 8'hec;
      17'd55885: data = 8'hef;
      17'd55886: data = 8'heb;
      17'd55887: data = 8'hef;
      17'd55888: data = 8'hec;
      17'd55889: data = 8'he7;
      17'd55890: data = 8'he4;
      17'd55891: data = 8'hef;
      17'd55892: data = 8'hf9;
      17'd55893: data = 8'h05;
      17'd55894: data = 8'h12;
      17'd55895: data = 8'h1f;
      17'd55896: data = 8'h2d;
      17'd55897: data = 8'h2c;
      17'd55898: data = 8'h2f;
      17'd55899: data = 8'h29;
      17'd55900: data = 8'h24;
      17'd55901: data = 8'h1c;
      17'd55902: data = 8'h0d;
      17'd55903: data = 8'h09;
      17'd55904: data = 8'h0c;
      17'd55905: data = 8'h0c;
      17'd55906: data = 8'h11;
      17'd55907: data = 8'h15;
      17'd55908: data = 8'h15;
      17'd55909: data = 8'h13;
      17'd55910: data = 8'h09;
      17'd55911: data = 8'h04;
      17'd55912: data = 8'h04;
      17'd55913: data = 8'h02;
      17'd55914: data = 8'hfc;
      17'd55915: data = 8'hf5;
      17'd55916: data = 8'hf1;
      17'd55917: data = 8'he7;
      17'd55918: data = 8'hd8;
      17'd55919: data = 8'hd2;
      17'd55920: data = 8'hd2;
      17'd55921: data = 8'hca;
      17'd55922: data = 8'hc4;
      17'd55923: data = 8'hc6;
      17'd55924: data = 8'hc9;
      17'd55925: data = 8'hcd;
      17'd55926: data = 8'hd3;
      17'd55927: data = 8'hd5;
      17'd55928: data = 8'hd5;
      17'd55929: data = 8'hd3;
      17'd55930: data = 8'hcb;
      17'd55931: data = 8'hc0;
      17'd55932: data = 8'hc0;
      17'd55933: data = 8'hc2;
      17'd55934: data = 8'hc6;
      17'd55935: data = 8'hcd;
      17'd55936: data = 8'hd8;
      17'd55937: data = 8'he0;
      17'd55938: data = 8'he4;
      17'd55939: data = 8'he9;
      17'd55940: data = 8'hf1;
      17'd55941: data = 8'hf9;
      17'd55942: data = 8'hf9;
      17'd55943: data = 8'hfd;
      17'd55944: data = 8'hfd;
      17'd55945: data = 8'hf5;
      17'd55946: data = 8'hfc;
      17'd55947: data = 8'hfe;
      17'd55948: data = 8'h00;
      17'd55949: data = 8'h09;
      17'd55950: data = 8'h05;
      17'd55951: data = 8'h05;
      17'd55952: data = 8'h06;
      17'd55953: data = 8'h09;
      17'd55954: data = 8'h0e;
      17'd55955: data = 8'h1a;
      17'd55956: data = 8'h22;
      17'd55957: data = 8'h27;
      17'd55958: data = 8'h1e;
      17'd55959: data = 8'h19;
      17'd55960: data = 8'h11;
      17'd55961: data = 8'h00;
      17'd55962: data = 8'h05;
      17'd55963: data = 8'h06;
      17'd55964: data = 8'h00;
      17'd55965: data = 8'hfc;
      17'd55966: data = 8'h01;
      17'd55967: data = 8'hfe;
      17'd55968: data = 8'h01;
      17'd55969: data = 8'h05;
      17'd55970: data = 8'h13;
      17'd55971: data = 8'h0c;
      17'd55972: data = 8'hfa;
      17'd55973: data = 8'h05;
      17'd55974: data = 8'hfe;
      17'd55975: data = 8'hde;
      17'd55976: data = 8'hec;
      17'd55977: data = 8'hf9;
      17'd55978: data = 8'hec;
      17'd55979: data = 8'hec;
      17'd55980: data = 8'heb;
      17'd55981: data = 8'hec;
      17'd55982: data = 8'hec;
      17'd55983: data = 8'hf1;
      17'd55984: data = 8'hf4;
      17'd55985: data = 8'hf9;
      17'd55986: data = 8'h01;
      17'd55987: data = 8'hed;
      17'd55988: data = 8'hfc;
      17'd55989: data = 8'h06;
      17'd55990: data = 8'hfc;
      17'd55991: data = 8'h12;
      17'd55992: data = 8'h0a;
      17'd55993: data = 8'h04;
      17'd55994: data = 8'h15;
      17'd55995: data = 8'h0a;
      17'd55996: data = 8'h1f;
      17'd55997: data = 8'h31;
      17'd55998: data = 8'h0a;
      17'd55999: data = 8'h19;
      17'd56000: data = 8'hfc;
      17'd56001: data = 8'hc5;
      17'd56002: data = 8'hef;
      17'd56003: data = 8'he5;
      17'd56004: data = 8'hed;
      17'd56005: data = 8'h1b;
      17'd56006: data = 8'h0a;
      17'd56007: data = 8'h1c;
      17'd56008: data = 8'h36;
      17'd56009: data = 8'h22;
      17'd56010: data = 8'h45;
      17'd56011: data = 8'h53;
      17'd56012: data = 8'h31;
      17'd56013: data = 8'h42;
      17'd56014: data = 8'h1a;
      17'd56015: data = 8'h01;
      17'd56016: data = 8'h12;
      17'd56017: data = 8'hfa;
      17'd56018: data = 8'h1a;
      17'd56019: data = 8'h1c;
      17'd56020: data = 8'h05;
      17'd56021: data = 8'h16;
      17'd56022: data = 8'h0a;
      17'd56023: data = 8'h01;
      17'd56024: data = 8'h27;
      17'd56025: data = 8'h36;
      17'd56026: data = 8'h39;
      17'd56027: data = 8'h3c;
      17'd56028: data = 8'h23;
      17'd56029: data = 8'h05;
      17'd56030: data = 8'hef;
      17'd56031: data = 8'he4;
      17'd56032: data = 8'he0;
      17'd56033: data = 8'hed;
      17'd56034: data = 8'hd6;
      17'd56035: data = 8'hd6;
      17'd56036: data = 8'hda;
      17'd56037: data = 8'hd5;
      17'd56038: data = 8'hf1;
      17'd56039: data = 8'hfa;
      17'd56040: data = 8'h02;
      17'd56041: data = 8'h00;
      17'd56042: data = 8'he7;
      17'd56043: data = 8'hd2;
      17'd56044: data = 8'hce;
      17'd56045: data = 8'hca;
      17'd56046: data = 8'hce;
      17'd56047: data = 8'he3;
      17'd56048: data = 8'hd5;
      17'd56049: data = 8'hce;
      17'd56050: data = 8'hcb;
      17'd56051: data = 8'hb9;
      17'd56052: data = 8'hc9;
      17'd56053: data = 8'he2;
      17'd56054: data = 8'hed;
      17'd56055: data = 8'h09;
      17'd56056: data = 8'h05;
      17'd56057: data = 8'h04;
      17'd56058: data = 8'h13;
      17'd56059: data = 8'h05;
      17'd56060: data = 8'h19;
      17'd56061: data = 8'h1a;
      17'd56062: data = 8'h11;
      17'd56063: data = 8'h0d;
      17'd56064: data = 8'h04;
      17'd56065: data = 8'h02;
      17'd56066: data = 8'h15;
      17'd56067: data = 8'h2b;
      17'd56068: data = 8'h3d;
      17'd56069: data = 8'h56;
      17'd56070: data = 8'h4f;
      17'd56071: data = 8'h47;
      17'd56072: data = 8'h42;
      17'd56073: data = 8'h35;
      17'd56074: data = 8'h3e;
      17'd56075: data = 8'h42;
      17'd56076: data = 8'h40;
      17'd56077: data = 8'h3c;
      17'd56078: data = 8'h2f;
      17'd56079: data = 8'h1f;
      17'd56080: data = 8'h1b;
      17'd56081: data = 8'h1a;
      17'd56082: data = 8'h1b;
      17'd56083: data = 8'h1f;
      17'd56084: data = 8'h1b;
      17'd56085: data = 8'h16;
      17'd56086: data = 8'h16;
      17'd56087: data = 8'h16;
      17'd56088: data = 8'h15;
      17'd56089: data = 8'h1a;
      17'd56090: data = 8'h12;
      17'd56091: data = 8'h05;
      17'd56092: data = 8'hf5;
      17'd56093: data = 8'hde;
      17'd56094: data = 8'hd6;
      17'd56095: data = 8'hd3;
      17'd56096: data = 8'hdb;
      17'd56097: data = 8'he4;
      17'd56098: data = 8'he9;
      17'd56099: data = 8'he9;
      17'd56100: data = 8'heb;
      17'd56101: data = 8'he9;
      17'd56102: data = 8'hec;
      17'd56103: data = 8'hf4;
      17'd56104: data = 8'hf4;
      17'd56105: data = 8'hf9;
      17'd56106: data = 8'hf5;
      17'd56107: data = 8'hef;
      17'd56108: data = 8'hf1;
      17'd56109: data = 8'hf1;
      17'd56110: data = 8'hf6;
      17'd56111: data = 8'hfd;
      17'd56112: data = 8'hfd;
      17'd56113: data = 8'h02;
      17'd56114: data = 8'h01;
      17'd56115: data = 8'h00;
      17'd56116: data = 8'h0c;
      17'd56117: data = 8'h16;
      17'd56118: data = 8'h23;
      17'd56119: data = 8'h2b;
      17'd56120: data = 8'h27;
      17'd56121: data = 8'h1e;
      17'd56122: data = 8'h13;
      17'd56123: data = 8'h0a;
      17'd56124: data = 8'h05;
      17'd56125: data = 8'h05;
      17'd56126: data = 8'h04;
      17'd56127: data = 8'h04;
      17'd56128: data = 8'h02;
      17'd56129: data = 8'h02;
      17'd56130: data = 8'h05;
      17'd56131: data = 8'h04;
      17'd56132: data = 8'h06;
      17'd56133: data = 8'h04;
      17'd56134: data = 8'hfa;
      17'd56135: data = 8'hf4;
      17'd56136: data = 8'hed;
      17'd56137: data = 8'he3;
      17'd56138: data = 8'he0;
      17'd56139: data = 8'he0;
      17'd56140: data = 8'hdb;
      17'd56141: data = 8'hd6;
      17'd56142: data = 8'hd1;
      17'd56143: data = 8'hcb;
      17'd56144: data = 8'hc9;
      17'd56145: data = 8'hca;
      17'd56146: data = 8'hd2;
      17'd56147: data = 8'hd8;
      17'd56148: data = 8'hdb;
      17'd56149: data = 8'hdb;
      17'd56150: data = 8'hdc;
      17'd56151: data = 8'hd5;
      17'd56152: data = 8'hd5;
      17'd56153: data = 8'hd5;
      17'd56154: data = 8'hd6;
      17'd56155: data = 8'hda;
      17'd56156: data = 8'hda;
      17'd56157: data = 8'hde;
      17'd56158: data = 8'hde;
      17'd56159: data = 8'he5;
      17'd56160: data = 8'hf4;
      17'd56161: data = 8'hfd;
      17'd56162: data = 8'hfe;
      17'd56163: data = 8'h05;
      17'd56164: data = 8'h00;
      17'd56165: data = 8'hfa;
      17'd56166: data = 8'hfa;
      17'd56167: data = 8'hfc;
      17'd56168: data = 8'hfe;
      17'd56169: data = 8'hfc;
      17'd56170: data = 8'hfe;
      17'd56171: data = 8'hfe;
      17'd56172: data = 8'hfc;
      17'd56173: data = 8'hf9;
      17'd56174: data = 8'h05;
      17'd56175: data = 8'h09;
      17'd56176: data = 8'h09;
      17'd56177: data = 8'h11;
      17'd56178: data = 8'h0d;
      17'd56179: data = 8'h0c;
      17'd56180: data = 8'h0a;
      17'd56181: data = 8'hfe;
      17'd56182: data = 8'h02;
      17'd56183: data = 8'h06;
      17'd56184: data = 8'hf5;
      17'd56185: data = 8'hf9;
      17'd56186: data = 8'hf5;
      17'd56187: data = 8'hed;
      17'd56188: data = 8'hf4;
      17'd56189: data = 8'hfd;
      17'd56190: data = 8'h04;
      17'd56191: data = 8'h00;
      17'd56192: data = 8'h00;
      17'd56193: data = 8'hfd;
      17'd56194: data = 8'hf5;
      17'd56195: data = 8'hf6;
      17'd56196: data = 8'hf5;
      17'd56197: data = 8'hfd;
      17'd56198: data = 8'h01;
      17'd56199: data = 8'he7;
      17'd56200: data = 8'hfc;
      17'd56201: data = 8'h00;
      17'd56202: data = 8'he2;
      17'd56203: data = 8'hfe;
      17'd56204: data = 8'hfe;
      17'd56205: data = 8'h00;
      17'd56206: data = 8'h05;
      17'd56207: data = 8'he2;
      17'd56208: data = 8'hfc;
      17'd56209: data = 8'hfd;
      17'd56210: data = 8'he9;
      17'd56211: data = 8'h1b;
      17'd56212: data = 8'h1c;
      17'd56213: data = 8'h06;
      17'd56214: data = 8'h2c;
      17'd56215: data = 8'h02;
      17'd56216: data = 8'hfd;
      17'd56217: data = 8'h13;
      17'd56218: data = 8'h0d;
      17'd56219: data = 8'h42;
      17'd56220: data = 8'h3c;
      17'd56221: data = 8'h24;
      17'd56222: data = 8'h2d;
      17'd56223: data = 8'he0;
      17'd56224: data = 8'hbb;
      17'd56225: data = 8'hbc;
      17'd56226: data = 8'hb0;
      17'd56227: data = 8'hd8;
      17'd56228: data = 8'hef;
      17'd56229: data = 8'hf4;
      17'd56230: data = 8'h22;
      17'd56231: data = 8'h22;
      17'd56232: data = 8'h26;
      17'd56233: data = 8'h47;
      17'd56234: data = 8'h4d;
      17'd56235: data = 8'h5a;
      17'd56236: data = 8'h31;
      17'd56237: data = 8'h0a;
      17'd56238: data = 8'hfd;
      17'd56239: data = 8'he2;
      17'd56240: data = 8'hdc;
      17'd56241: data = 8'hfa;
      17'd56242: data = 8'h11;
      17'd56243: data = 8'h16;
      17'd56244: data = 8'h06;
      17'd56245: data = 8'h01;
      17'd56246: data = 8'hfc;
      17'd56247: data = 8'h0d;
      17'd56248: data = 8'h33;
      17'd56249: data = 8'h4b;
      17'd56250: data = 8'h5c;
      17'd56251: data = 8'h4b;
      17'd56252: data = 8'h26;
      17'd56253: data = 8'hf9;
      17'd56254: data = 8'hd6;
      17'd56255: data = 8'hd8;
      17'd56256: data = 8'hde;
      17'd56257: data = 8'hce;
      17'd56258: data = 8'hd5;
      17'd56259: data = 8'hd3;
      17'd56260: data = 8'hc0;
      17'd56261: data = 8'hd5;
      17'd56262: data = 8'hed;
      17'd56263: data = 8'h11;
      17'd56264: data = 8'h24;
      17'd56265: data = 8'h0c;
      17'd56266: data = 8'hfd;
      17'd56267: data = 8'he2;
      17'd56268: data = 8'hb9;
      17'd56269: data = 8'hbd;
      17'd56270: data = 8'hc2;
      17'd56271: data = 8'hd1;
      17'd56272: data = 8'hd2;
      17'd56273: data = 8'hb4;
      17'd56274: data = 8'hb0;
      17'd56275: data = 8'haa;
      17'd56276: data = 8'hb0;
      17'd56277: data = 8'hd2;
      17'd56278: data = 8'hf6;
      17'd56279: data = 8'h0e;
      17'd56280: data = 8'h1b;
      17'd56281: data = 8'h16;
      17'd56282: data = 8'h12;
      17'd56283: data = 8'h13;
      17'd56284: data = 8'h13;
      17'd56285: data = 8'h15;
      17'd56286: data = 8'h11;
      17'd56287: data = 8'h05;
      17'd56288: data = 8'hfa;
      17'd56289: data = 8'hef;
      17'd56290: data = 8'hf6;
      17'd56291: data = 8'h13;
      17'd56292: data = 8'h3a;
      17'd56293: data = 8'h53;
      17'd56294: data = 8'h5c;
      17'd56295: data = 8'h5d;
      17'd56296: data = 8'h4f;
      17'd56297: data = 8'h45;
      17'd56298: data = 8'h3e;
      17'd56299: data = 8'h42;
      17'd56300: data = 8'h45;
      17'd56301: data = 8'h3a;
      17'd56302: data = 8'h27;
      17'd56303: data = 8'h1e;
      17'd56304: data = 8'h04;
      17'd56305: data = 8'hfd;
      17'd56306: data = 8'h04;
      17'd56307: data = 8'h09;
      17'd56308: data = 8'h16;
      17'd56309: data = 8'h16;
      17'd56310: data = 8'h15;
      17'd56311: data = 8'h19;
      17'd56312: data = 8'h16;
      17'd56313: data = 8'h15;
      17'd56314: data = 8'h19;
      17'd56315: data = 8'h0d;
      17'd56316: data = 8'hfe;
      17'd56317: data = 8'heb;
      17'd56318: data = 8'hce;
      17'd56319: data = 8'hc5;
      17'd56320: data = 8'hc6;
      17'd56321: data = 8'hd1;
      17'd56322: data = 8'hdb;
      17'd56323: data = 8'he3;
      17'd56324: data = 8'hed;
      17'd56325: data = 8'hf2;
      17'd56326: data = 8'hef;
      17'd56327: data = 8'hfc;
      17'd56328: data = 8'h0a;
      17'd56329: data = 8'h11;
      17'd56330: data = 8'h13;
      17'd56331: data = 8'h12;
      17'd56332: data = 8'h05;
      17'd56333: data = 8'hfc;
      17'd56334: data = 8'hf6;
      17'd56335: data = 8'hf1;
      17'd56336: data = 8'hf9;
      17'd56337: data = 8'h01;
      17'd56338: data = 8'h01;
      17'd56339: data = 8'h02;
      17'd56340: data = 8'h09;
      17'd56341: data = 8'h16;
      17'd56342: data = 8'h23;
      17'd56343: data = 8'h2c;
      17'd56344: data = 8'h35;
      17'd56345: data = 8'h31;
      17'd56346: data = 8'h23;
      17'd56347: data = 8'h13;
      17'd56348: data = 8'h09;
      17'd56349: data = 8'h01;
      17'd56350: data = 8'hfc;
      17'd56351: data = 8'hfa;
      17'd56352: data = 8'hf9;
      17'd56353: data = 8'hf2;
      17'd56354: data = 8'hed;
      17'd56355: data = 8'hed;
      17'd56356: data = 8'hf1;
      17'd56357: data = 8'hf9;
      17'd56358: data = 8'hfd;
      17'd56359: data = 8'hfa;
      17'd56360: data = 8'hf5;
      17'd56361: data = 8'hec;
      17'd56362: data = 8'hde;
      17'd56363: data = 8'hda;
      17'd56364: data = 8'hd2;
      17'd56365: data = 8'hd1;
      17'd56366: data = 8'hcb;
      17'd56367: data = 8'hc2;
      17'd56368: data = 8'hc5;
      17'd56369: data = 8'hc1;
      17'd56370: data = 8'hcb;
      17'd56371: data = 8'hd6;
      17'd56372: data = 8'hdc;
      17'd56373: data = 8'he9;
      17'd56374: data = 8'hec;
      17'd56375: data = 8'he4;
      17'd56376: data = 8'he4;
      17'd56377: data = 8'he3;
      17'd56378: data = 8'he4;
      17'd56379: data = 8'he5;
      17'd56380: data = 8'he4;
      17'd56381: data = 8'he5;
      17'd56382: data = 8'he5;
      17'd56383: data = 8'he7;
      17'd56384: data = 8'hf1;
      17'd56385: data = 8'h00;
      17'd56386: data = 8'h05;
      17'd56387: data = 8'h0a;
      17'd56388: data = 8'h0a;
      17'd56389: data = 8'h02;
      17'd56390: data = 8'hfd;
      17'd56391: data = 8'hfd;
      17'd56392: data = 8'hfc;
      17'd56393: data = 8'h00;
      17'd56394: data = 8'h02;
      17'd56395: data = 8'hfd;
      17'd56396: data = 8'hf9;
      17'd56397: data = 8'hf6;
      17'd56398: data = 8'hf6;
      17'd56399: data = 8'hfd;
      17'd56400: data = 8'hfe;
      17'd56401: data = 8'h13;
      17'd56402: data = 8'h0c;
      17'd56403: data = 8'h02;
      17'd56404: data = 8'h19;
      17'd56405: data = 8'hfa;
      17'd56406: data = 8'hf6;
      17'd56407: data = 8'h0c;
      17'd56408: data = 8'hf6;
      17'd56409: data = 8'hf9;
      17'd56410: data = 8'hf9;
      17'd56411: data = 8'he3;
      17'd56412: data = 8'hf9;
      17'd56413: data = 8'heb;
      17'd56414: data = 8'hf4;
      17'd56415: data = 8'h1b;
      17'd56416: data = 8'hfd;
      17'd56417: data = 8'h04;
      17'd56418: data = 8'h1b;
      17'd56419: data = 8'he5;
      17'd56420: data = 8'h06;
      17'd56421: data = 8'h0c;
      17'd56422: data = 8'he3;
      17'd56423: data = 8'h1f;
      17'd56424: data = 8'hf2;
      17'd56425: data = 8'hf1;
      17'd56426: data = 8'h0a;
      17'd56427: data = 8'he4;
      17'd56428: data = 8'h0c;
      17'd56429: data = 8'h0c;
      17'd56430: data = 8'hf5;
      17'd56431: data = 8'h1f;
      17'd56432: data = 8'h0a;
      17'd56433: data = 8'hfa;
      17'd56434: data = 8'h0e;
      17'd56435: data = 8'h0e;
      17'd56436: data = 8'h13;
      17'd56437: data = 8'h0c;
      17'd56438: data = 8'h13;
      17'd56439: data = 8'h1e;
      17'd56440: data = 8'h19;
      17'd56441: data = 8'h09;
      17'd56442: data = 8'h0d;
      17'd56443: data = 8'h02;
      17'd56444: data = 8'he0;
      17'd56445: data = 8'hde;
      17'd56446: data = 8'hcd;
      17'd56447: data = 8'hd5;
      17'd56448: data = 8'he4;
      17'd56449: data = 8'he5;
      17'd56450: data = 8'hfe;
      17'd56451: data = 8'h0c;
      17'd56452: data = 8'h23;
      17'd56453: data = 8'h1f;
      17'd56454: data = 8'h31;
      17'd56455: data = 8'h3e;
      17'd56456: data = 8'h2d;
      17'd56457: data = 8'h27;
      17'd56458: data = 8'h09;
      17'd56459: data = 8'h11;
      17'd56460: data = 8'hfc;
      17'd56461: data = 8'hf2;
      17'd56462: data = 8'h0d;
      17'd56463: data = 8'h05;
      17'd56464: data = 8'h0e;
      17'd56465: data = 8'h13;
      17'd56466: data = 8'h02;
      17'd56467: data = 8'h19;
      17'd56468: data = 8'h1e;
      17'd56469: data = 8'h2c;
      17'd56470: data = 8'h34;
      17'd56471: data = 8'h3a;
      17'd56472: data = 8'h36;
      17'd56473: data = 8'h11;
      17'd56474: data = 8'h09;
      17'd56475: data = 8'hf2;
      17'd56476: data = 8'hf9;
      17'd56477: data = 8'he2;
      17'd56478: data = 8'hd8;
      17'd56479: data = 8'hdc;
      17'd56480: data = 8'hc9;
      17'd56481: data = 8'hd3;
      17'd56482: data = 8'hda;
      17'd56483: data = 8'hf1;
      17'd56484: data = 8'h06;
      17'd56485: data = 8'h00;
      17'd56486: data = 8'h00;
      17'd56487: data = 8'hf2;
      17'd56488: data = 8'hdc;
      17'd56489: data = 8'hd3;
      17'd56490: data = 8'hc4;
      17'd56491: data = 8'hd1;
      17'd56492: data = 8'hc6;
      17'd56493: data = 8'hca;
      17'd56494: data = 8'hc1;
      17'd56495: data = 8'hb4;
      17'd56496: data = 8'hc1;
      17'd56497: data = 8'hc1;
      17'd56498: data = 8'hdc;
      17'd56499: data = 8'he7;
      17'd56500: data = 8'hfc;
      17'd56501: data = 8'h0d;
      17'd56502: data = 8'h04;
      17'd56503: data = 8'h0d;
      17'd56504: data = 8'h12;
      17'd56505: data = 8'h16;
      17'd56506: data = 8'h19;
      17'd56507: data = 8'h12;
      17'd56508: data = 8'h0e;
      17'd56509: data = 8'h01;
      17'd56510: data = 8'hfa;
      17'd56511: data = 8'hfd;
      17'd56512: data = 8'h0e;
      17'd56513: data = 8'h26;
      17'd56514: data = 8'h34;
      17'd56515: data = 8'h45;
      17'd56516: data = 8'h42;
      17'd56517: data = 8'h45;
      17'd56518: data = 8'h42;
      17'd56519: data = 8'h35;
      17'd56520: data = 8'h3e;
      17'd56521: data = 8'h34;
      17'd56522: data = 8'h2d;
      17'd56523: data = 8'h23;
      17'd56524: data = 8'h15;
      17'd56525: data = 8'h0c;
      17'd56526: data = 8'h04;
      17'd56527: data = 8'h05;
      17'd56528: data = 8'h05;
      17'd56529: data = 8'h0a;
      17'd56530: data = 8'h06;
      17'd56531: data = 8'h06;
      17'd56532: data = 8'h05;
      17'd56533: data = 8'h0a;
      17'd56534: data = 8'h11;
      17'd56535: data = 8'h0a;
      17'd56536: data = 8'h0a;
      17'd56537: data = 8'h0a;
      17'd56538: data = 8'hf5;
      17'd56539: data = 8'he7;
      17'd56540: data = 8'he0;
      17'd56541: data = 8'hd6;
      17'd56542: data = 8'hdc;
      17'd56543: data = 8'he0;
      17'd56544: data = 8'hed;
      17'd56545: data = 8'hf4;
      17'd56546: data = 8'hf6;
      17'd56547: data = 8'hfa;
      17'd56548: data = 8'hfe;
      17'd56549: data = 8'h09;
      17'd56550: data = 8'h0e;
      17'd56551: data = 8'h15;
      17'd56552: data = 8'h11;
      17'd56553: data = 8'h13;
      17'd56554: data = 8'h0e;
      17'd56555: data = 8'h04;
      17'd56556: data = 8'h0c;
      17'd56557: data = 8'h0c;
      17'd56558: data = 8'h0e;
      17'd56559: data = 8'h0e;
      17'd56560: data = 8'h0e;
      17'd56561: data = 8'h0d;
      17'd56562: data = 8'h0d;
      17'd56563: data = 8'h16;
      17'd56564: data = 8'h1b;
      17'd56565: data = 8'h1a;
      17'd56566: data = 8'h15;
      17'd56567: data = 8'h1a;
      17'd56568: data = 8'h0e;
      17'd56569: data = 8'h00;
      17'd56570: data = 8'h0d;
      17'd56571: data = 8'h0c;
      17'd56572: data = 8'hfe;
      17'd56573: data = 8'h05;
      17'd56574: data = 8'hfe;
      17'd56575: data = 8'hf9;
      17'd56576: data = 8'hf2;
      17'd56577: data = 8'heb;
      17'd56578: data = 8'he9;
      17'd56579: data = 8'he7;
      17'd56580: data = 8'hec;
      17'd56581: data = 8'heb;
      17'd56582: data = 8'he7;
      17'd56583: data = 8'he2;
      17'd56584: data = 8'he2;
      17'd56585: data = 8'hde;
      17'd56586: data = 8'hda;
      17'd56587: data = 8'he0;
      17'd56588: data = 8'hdb;
      17'd56589: data = 8'hd5;
      17'd56590: data = 8'hd6;
      17'd56591: data = 8'hd3;
      17'd56592: data = 8'hd5;
      17'd56593: data = 8'hda;
      17'd56594: data = 8'hde;
      17'd56595: data = 8'he3;
      17'd56596: data = 8'he4;
      17'd56597: data = 8'he0;
      17'd56598: data = 8'he2;
      17'd56599: data = 8'heb;
      17'd56600: data = 8'he9;
      17'd56601: data = 8'hf2;
      17'd56602: data = 8'hf6;
      17'd56603: data = 8'hfa;
      17'd56604: data = 8'hfc;
      17'd56605: data = 8'hfa;
      17'd56606: data = 8'hfd;
      17'd56607: data = 8'hf9;
      17'd56608: data = 8'hf9;
      17'd56609: data = 8'hfa;
      17'd56610: data = 8'hf5;
      17'd56611: data = 8'hfa;
      17'd56612: data = 8'hf9;
      17'd56613: data = 8'hf9;
      17'd56614: data = 8'hf6;
      17'd56615: data = 8'hf9;
      17'd56616: data = 8'h01;
      17'd56617: data = 8'hf4;
      17'd56618: data = 8'hfa;
      17'd56619: data = 8'h02;
      17'd56620: data = 8'hf9;
      17'd56621: data = 8'hf9;
      17'd56622: data = 8'hfe;
      17'd56623: data = 8'hfe;
      17'd56624: data = 8'hfc;
      17'd56625: data = 8'hfe;
      17'd56626: data = 8'hfc;
      17'd56627: data = 8'hf9;
      17'd56628: data = 8'hfd;
      17'd56629: data = 8'hef;
      17'd56630: data = 8'hfa;
      17'd56631: data = 8'hfe;
      17'd56632: data = 8'hf5;
      17'd56633: data = 8'h06;
      17'd56634: data = 8'hf9;
      17'd56635: data = 8'h09;
      17'd56636: data = 8'h0d;
      17'd56637: data = 8'hf9;
      17'd56638: data = 8'h0e;
      17'd56639: data = 8'h05;
      17'd56640: data = 8'h09;
      17'd56641: data = 8'h11;
      17'd56642: data = 8'hfe;
      17'd56643: data = 8'h0e;
      17'd56644: data = 8'h05;
      17'd56645: data = 8'hfe;
      17'd56646: data = 8'h13;
      17'd56647: data = 8'h02;
      17'd56648: data = 8'h1a;
      17'd56649: data = 8'h0c;
      17'd56650: data = 8'h06;
      17'd56651: data = 8'h24;
      17'd56652: data = 8'hf6;
      17'd56653: data = 8'hf4;
      17'd56654: data = 8'h29;
      17'd56655: data = 8'hf6;
      17'd56656: data = 8'hfc;
      17'd56657: data = 8'h27;
      17'd56658: data = 8'h0e;
      17'd56659: data = 8'h19;
      17'd56660: data = 8'h2f;
      17'd56661: data = 8'h2f;
      17'd56662: data = 8'h4d;
      17'd56663: data = 8'h2d;
      17'd56664: data = 8'h27;
      17'd56665: data = 8'h1e;
      17'd56666: data = 8'hcb;
      17'd56667: data = 8'hc6;
      17'd56668: data = 8'hbc;
      17'd56669: data = 8'h9d;
      17'd56670: data = 8'hbd;
      17'd56671: data = 8'he0;
      17'd56672: data = 8'hed;
      17'd56673: data = 8'h05;
      17'd56674: data = 8'h24;
      17'd56675: data = 8'h33;
      17'd56676: data = 8'h29;
      17'd56677: data = 8'h33;
      17'd56678: data = 8'h2c;
      17'd56679: data = 8'h23;
      17'd56680: data = 8'h12;
      17'd56681: data = 8'h00;
      17'd56682: data = 8'h04;
      17'd56683: data = 8'hf6;
      17'd56684: data = 8'hfe;
      17'd56685: data = 8'h02;
      17'd56686: data = 8'hfc;
      17'd56687: data = 8'h06;
      17'd56688: data = 8'h02;
      17'd56689: data = 8'hfd;
      17'd56690: data = 8'h19;
      17'd56691: data = 8'h2d;
      17'd56692: data = 8'h33;
      17'd56693: data = 8'h4d;
      17'd56694: data = 8'h4d;
      17'd56695: data = 8'h39;
      17'd56696: data = 8'h26;
      17'd56697: data = 8'h02;
      17'd56698: data = 8'hec;
      17'd56699: data = 8'hda;
      17'd56700: data = 8'hc5;
      17'd56701: data = 8'hce;
      17'd56702: data = 8'hc6;
      17'd56703: data = 8'hd3;
      17'd56704: data = 8'he2;
      17'd56705: data = 8'he3;
      17'd56706: data = 8'hfd;
      17'd56707: data = 8'h01;
      17'd56708: data = 8'h02;
      17'd56709: data = 8'hfe;
      17'd56710: data = 8'hf2;
      17'd56711: data = 8'he2;
      17'd56712: data = 8'hd1;
      17'd56713: data = 8'hd3;
      17'd56714: data = 8'hc5;
      17'd56715: data = 8'hc1;
      17'd56716: data = 8'hc4;
      17'd56717: data = 8'hbb;
      17'd56718: data = 8'hb0;
      17'd56719: data = 8'hb3;
      17'd56720: data = 8'hc4;
      17'd56721: data = 8'hd1;
      17'd56722: data = 8'hde;
      17'd56723: data = 8'h06;
      17'd56724: data = 8'h16;
      17'd56725: data = 8'h13;
      17'd56726: data = 8'h26;
      17'd56727: data = 8'h27;
      17'd56728: data = 8'h13;
      17'd56729: data = 8'h0c;
      17'd56730: data = 8'h0c;
      17'd56731: data = 8'hfd;
      17'd56732: data = 8'hf4;
      17'd56733: data = 8'hf6;
      17'd56734: data = 8'h05;
      17'd56735: data = 8'h11;
      17'd56736: data = 8'h22;
      17'd56737: data = 8'h40;
      17'd56738: data = 8'h42;
      17'd56739: data = 8'h43;
      17'd56740: data = 8'h4b;
      17'd56741: data = 8'h43;
      17'd56742: data = 8'h3e;
      17'd56743: data = 8'h3c;
      17'd56744: data = 8'h35;
      17'd56745: data = 8'h2d;
      17'd56746: data = 8'h22;
      17'd56747: data = 8'h13;
      17'd56748: data = 8'h0a;
      17'd56749: data = 8'h01;
      17'd56750: data = 8'hf2;
      17'd56751: data = 8'hf2;
      17'd56752: data = 8'hf9;
      17'd56753: data = 8'hfa;
      17'd56754: data = 8'h00;
      17'd56755: data = 8'h0a;
      17'd56756: data = 8'h1a;
      17'd56757: data = 8'h1b;
      17'd56758: data = 8'h0e;
      17'd56759: data = 8'h16;
      17'd56760: data = 8'h09;
      17'd56761: data = 8'hef;
      17'd56762: data = 8'he5;
      17'd56763: data = 8'hde;
      17'd56764: data = 8'hd1;
      17'd56765: data = 8'hd2;
      17'd56766: data = 8'hde;
      17'd56767: data = 8'he4;
      17'd56768: data = 8'heb;
      17'd56769: data = 8'hf9;
      17'd56770: data = 8'h09;
      17'd56771: data = 8'h0c;
      17'd56772: data = 8'h13;
      17'd56773: data = 8'h23;
      17'd56774: data = 8'h1c;
      17'd56775: data = 8'h13;
      17'd56776: data = 8'h19;
      17'd56777: data = 8'h12;
      17'd56778: data = 8'h0a;
      17'd56779: data = 8'h0a;
      17'd56780: data = 8'h09;
      17'd56781: data = 8'h02;
      17'd56782: data = 8'h01;
      17'd56783: data = 8'h02;
      17'd56784: data = 8'h01;
      17'd56785: data = 8'h0d;
      17'd56786: data = 8'h1a;
      17'd56787: data = 8'h1b;
      17'd56788: data = 8'h2c;
      17'd56789: data = 8'h31;
      17'd56790: data = 8'h26;
      17'd56791: data = 8'h1c;
      17'd56792: data = 8'h13;
      17'd56793: data = 8'h09;
      17'd56794: data = 8'hf4;
      17'd56795: data = 8'hf2;
      17'd56796: data = 8'hf2;
      17'd56797: data = 8'he5;
      17'd56798: data = 8'he7;
      17'd56799: data = 8'hf1;
      17'd56800: data = 8'hef;
      17'd56801: data = 8'hec;
      17'd56802: data = 8'hf4;
      17'd56803: data = 8'hf6;
      17'd56804: data = 8'hef;
      17'd56805: data = 8'hf1;
      17'd56806: data = 8'hed;
      17'd56807: data = 8'he3;
      17'd56808: data = 8'hde;
      17'd56809: data = 8'hd8;
      17'd56810: data = 8'hd8;
      17'd56811: data = 8'hd3;
      17'd56812: data = 8'hd1;
      17'd56813: data = 8'hd3;
      17'd56814: data = 8'hd1;
      17'd56815: data = 8'hd6;
      17'd56816: data = 8'he0;
      17'd56817: data = 8'he3;
      17'd56818: data = 8'hec;
      17'd56819: data = 8'hf4;
      17'd56820: data = 8'hf5;
      17'd56821: data = 8'hfc;
      17'd56822: data = 8'hf6;
      17'd56823: data = 8'hef;
      17'd56824: data = 8'hef;
      17'd56825: data = 8'hef;
      17'd56826: data = 8'hed;
      17'd56827: data = 8'hf1;
      17'd56828: data = 8'hf9;
      17'd56829: data = 8'hfc;
      17'd56830: data = 8'hfd;
      17'd56831: data = 8'hfd;
      17'd56832: data = 8'h01;
      17'd56833: data = 8'hfe;
      17'd56834: data = 8'hfc;
      17'd56835: data = 8'h01;
      17'd56836: data = 8'hfe;
      17'd56837: data = 8'hf5;
      17'd56838: data = 8'hf6;
      17'd56839: data = 8'hf6;
      17'd56840: data = 8'hed;
      17'd56841: data = 8'hf1;
      17'd56842: data = 8'hf5;
      17'd56843: data = 8'hf5;
      17'd56844: data = 8'hf9;
      17'd56845: data = 8'hfc;
      17'd56846: data = 8'hfe;
      17'd56847: data = 8'hfd;
      17'd56848: data = 8'h01;
      17'd56849: data = 8'h04;
      17'd56850: data = 8'h00;
      17'd56851: data = 8'h00;
      17'd56852: data = 8'hfd;
      17'd56853: data = 8'hf4;
      17'd56854: data = 8'hf9;
      17'd56855: data = 8'hf4;
      17'd56856: data = 8'hed;
      17'd56857: data = 8'h06;
      17'd56858: data = 8'hfd;
      17'd56859: data = 8'hfd;
      17'd56860: data = 8'h12;
      17'd56861: data = 8'h0c;
      17'd56862: data = 8'h11;
      17'd56863: data = 8'h09;
      17'd56864: data = 8'h19;
      17'd56865: data = 8'h11;
      17'd56866: data = 8'hfd;
      17'd56867: data = 8'h15;
      17'd56868: data = 8'hf9;
      17'd56869: data = 8'hfd;
      17'd56870: data = 8'h09;
      17'd56871: data = 8'hf2;
      17'd56872: data = 8'h06;
      17'd56873: data = 8'h0a;
      17'd56874: data = 8'hfc;
      17'd56875: data = 8'h0d;
      17'd56876: data = 8'h0a;
      17'd56877: data = 8'h1a;
      17'd56878: data = 8'h0c;
      17'd56879: data = 8'h23;
      17'd56880: data = 8'h3a;
      17'd56881: data = 8'h15;
      17'd56882: data = 8'h40;
      17'd56883: data = 8'h42;
      17'd56884: data = 8'h0c;
      17'd56885: data = 8'h19;
      17'd56886: data = 8'hef;
      17'd56887: data = 8'hd3;
      17'd56888: data = 8'hbb;
      17'd56889: data = 8'ha8;
      17'd56890: data = 8'hce;
      17'd56891: data = 8'hc5;
      17'd56892: data = 8'hdb;
      17'd56893: data = 8'h29;
      17'd56894: data = 8'h1c;
      17'd56895: data = 8'h33;
      17'd56896: data = 8'h53;
      17'd56897: data = 8'h2f;
      17'd56898: data = 8'h2f;
      17'd56899: data = 8'h1f;
      17'd56900: data = 8'h12;
      17'd56901: data = 8'h12;
      17'd56902: data = 8'hf5;
      17'd56903: data = 8'h05;
      17'd56904: data = 8'h01;
      17'd56905: data = 8'hf1;
      17'd56906: data = 8'h04;
      17'd56907: data = 8'hfe;
      17'd56908: data = 8'h0a;
      17'd56909: data = 8'h19;
      17'd56910: data = 8'h1c;
      17'd56911: data = 8'h36;
      17'd56912: data = 8'h3d;
      17'd56913: data = 8'h3c;
      17'd56914: data = 8'h34;
      17'd56915: data = 8'h36;
      17'd56916: data = 8'h1f;
      17'd56917: data = 8'hfd;
      17'd56918: data = 8'hf4;
      17'd56919: data = 8'hda;
      17'd56920: data = 8'hc1;
      17'd56921: data = 8'hc0;
      17'd56922: data = 8'hcb;
      17'd56923: data = 8'hdb;
      17'd56924: data = 8'hde;
      17'd56925: data = 8'hf9;
      17'd56926: data = 8'h0c;
      17'd56927: data = 8'hfe;
      17'd56928: data = 8'h04;
      17'd56929: data = 8'h02;
      17'd56930: data = 8'he9;
      17'd56931: data = 8'he3;
      17'd56932: data = 8'hd8;
      17'd56933: data = 8'hca;
      17'd56934: data = 8'hc9;
      17'd56935: data = 8'hbb;
      17'd56936: data = 8'hb9;
      17'd56937: data = 8'hb9;
      17'd56938: data = 8'hb3;
      17'd56939: data = 8'hc5;
      17'd56940: data = 8'hca;
      17'd56941: data = 8'hd5;
      17'd56942: data = 8'hef;
      17'd56943: data = 8'hf2;
      17'd56944: data = 8'h09;
      17'd56945: data = 8'h13;
      17'd56946: data = 8'h0d;
      17'd56947: data = 8'h15;
      17'd56948: data = 8'h0d;
      17'd56949: data = 8'h00;
      17'd56950: data = 8'hf4;
      17'd56951: data = 8'hf4;
      17'd56952: data = 8'hf6;
      17'd56953: data = 8'hf1;
      17'd56954: data = 8'hfe;
      17'd56955: data = 8'h19;
      17'd56956: data = 8'h27;
      17'd56957: data = 8'h31;
      17'd56958: data = 8'h3e;
      17'd56959: data = 8'h4b;
      17'd56960: data = 8'h40;
      17'd56961: data = 8'h3e;
      17'd56962: data = 8'h40;
      17'd56963: data = 8'h31;
      17'd56964: data = 8'h27;
      17'd56965: data = 8'h1f;
      17'd56966: data = 8'h19;
      17'd56967: data = 8'h11;
      17'd56968: data = 8'h09;
      17'd56969: data = 8'h06;
      17'd56970: data = 8'h05;
      17'd56971: data = 8'h01;
      17'd56972: data = 8'h05;
      17'd56973: data = 8'h0a;
      17'd56974: data = 8'h0d;
      17'd56975: data = 8'h12;
      17'd56976: data = 8'h16;
      17'd56977: data = 8'h19;
      17'd56978: data = 8'h15;
      17'd56979: data = 8'h05;
      17'd56980: data = 8'hfd;
      17'd56981: data = 8'hf6;
      17'd56982: data = 8'he2;
      17'd56983: data = 8'hd6;
      17'd56984: data = 8'hd6;
      17'd56985: data = 8'hda;
      17'd56986: data = 8'hd8;
      17'd56987: data = 8'he2;
      17'd56988: data = 8'hf4;
      17'd56989: data = 8'hfa;
      17'd56990: data = 8'h00;
      17'd56991: data = 8'h09;
      17'd56992: data = 8'h0e;
      17'd56993: data = 8'h0c;
      17'd56994: data = 8'h09;
      17'd56995: data = 8'h0e;
      17'd56996: data = 8'h06;
      17'd56997: data = 8'hfd;
      17'd56998: data = 8'h04;
      17'd56999: data = 8'h01;
      17'd57000: data = 8'h00;
      17'd57001: data = 8'h05;
      17'd57002: data = 8'h04;
      17'd57003: data = 8'h06;
      17'd57004: data = 8'h0a;
      17'd57005: data = 8'h0e;
      17'd57006: data = 8'h1c;
      17'd57007: data = 8'h1e;
      17'd57008: data = 8'h1f;
      17'd57009: data = 8'h24;
      17'd57010: data = 8'h1f;
      17'd57011: data = 8'h16;
      17'd57012: data = 8'h11;
      17'd57013: data = 8'h09;
      17'd57014: data = 8'h02;
      17'd57015: data = 8'hf9;
      17'd57016: data = 8'hf5;
      17'd57017: data = 8'hf9;
      17'd57018: data = 8'hf1;
      17'd57019: data = 8'hf2;
      17'd57020: data = 8'hfa;
      17'd57021: data = 8'hfa;
      17'd57022: data = 8'hfd;
      17'd57023: data = 8'hfe;
      17'd57024: data = 8'hf6;
      17'd57025: data = 8'hf1;
      17'd57026: data = 8'he7;
      17'd57027: data = 8'he2;
      17'd57028: data = 8'hde;
      17'd57029: data = 8'hdb;
      17'd57030: data = 8'hda;
      17'd57031: data = 8'hd8;
      17'd57032: data = 8'hd5;
      17'd57033: data = 8'hd6;
      17'd57034: data = 8'hd5;
      17'd57035: data = 8'hd6;
      17'd57036: data = 8'he2;
      17'd57037: data = 8'he3;
      17'd57038: data = 8'he5;
      17'd57039: data = 8'heb;
      17'd57040: data = 8'he7;
      17'd57041: data = 8'he7;
      17'd57042: data = 8'he7;
      17'd57043: data = 8'he3;
      17'd57044: data = 8'he4;
      17'd57045: data = 8'he9;
      17'd57046: data = 8'heb;
      17'd57047: data = 8'hec;
      17'd57048: data = 8'hf1;
      17'd57049: data = 8'hf6;
      17'd57050: data = 8'hfc;
      17'd57051: data = 8'hfd;
      17'd57052: data = 8'hfe;
      17'd57053: data = 8'h00;
      17'd57054: data = 8'hfc;
      17'd57055: data = 8'hf9;
      17'd57056: data = 8'hf4;
      17'd57057: data = 8'hf1;
      17'd57058: data = 8'hf2;
      17'd57059: data = 8'hf1;
      17'd57060: data = 8'hf2;
      17'd57061: data = 8'hf9;
      17'd57062: data = 8'hf6;
      17'd57063: data = 8'hf9;
      17'd57064: data = 8'hfd;
      17'd57065: data = 8'hfe;
      17'd57066: data = 8'h02;
      17'd57067: data = 8'h06;
      17'd57068: data = 8'h05;
      17'd57069: data = 8'h06;
      17'd57070: data = 8'h02;
      17'd57071: data = 8'hfe;
      17'd57072: data = 8'hfd;
      17'd57073: data = 8'hfd;
      17'd57074: data = 8'hf6;
      17'd57075: data = 8'hfd;
      17'd57076: data = 8'hfe;
      17'd57077: data = 8'h00;
      17'd57078: data = 8'h0c;
      17'd57079: data = 8'h09;
      17'd57080: data = 8'h11;
      17'd57081: data = 8'h15;
      17'd57082: data = 8'h0e;
      17'd57083: data = 8'h15;
      17'd57084: data = 8'h13;
      17'd57085: data = 8'hfc;
      17'd57086: data = 8'h19;
      17'd57087: data = 8'hfe;
      17'd57088: data = 8'hfc;
      17'd57089: data = 8'h22;
      17'd57090: data = 8'hf9;
      17'd57091: data = 8'h0d;
      17'd57092: data = 8'h22;
      17'd57093: data = 8'hf6;
      17'd57094: data = 8'h1c;
      17'd57095: data = 8'h0c;
      17'd57096: data = 8'hfa;
      17'd57097: data = 8'h2b;
      17'd57098: data = 8'hf6;
      17'd57099: data = 8'h04;
      17'd57100: data = 8'h3a;
      17'd57101: data = 8'he5;
      17'd57102: data = 8'h1a;
      17'd57103: data = 8'h1c;
      17'd57104: data = 8'he0;
      17'd57105: data = 8'h1c;
      17'd57106: data = 8'hec;
      17'd57107: data = 8'hed;
      17'd57108: data = 8'h12;
      17'd57109: data = 8'hd3;
      17'd57110: data = 8'h06;
      17'd57111: data = 8'h2b;
      17'd57112: data = 8'hd6;
      17'd57113: data = 8'h22;
      17'd57114: data = 8'h06;
      17'd57115: data = 8'hc4;
      17'd57116: data = 8'h0c;
      17'd57117: data = 8'he5;
      17'd57118: data = 8'hf9;
      17'd57119: data = 8'h24;
      17'd57120: data = 8'h06;
      17'd57121: data = 8'h3c;
      17'd57122: data = 8'h2b;
      17'd57123: data = 8'hfc;
      17'd57124: data = 8'h35;
      17'd57125: data = 8'h11;
      17'd57126: data = 8'he4;
      17'd57127: data = 8'h2f;
      17'd57128: data = 8'h0d;
      17'd57129: data = 8'h02;
      17'd57130: data = 8'h2d;
      17'd57131: data = 8'h0a;
      17'd57132: data = 8'h1e;
      17'd57133: data = 8'h1f;
      17'd57134: data = 8'h04;
      17'd57135: data = 8'h2b;
      17'd57136: data = 8'h15;
      17'd57137: data = 8'hf5;
      17'd57138: data = 8'h31;
      17'd57139: data = 8'hfe;
      17'd57140: data = 8'h01;
      17'd57141: data = 8'h29;
      17'd57142: data = 8'hef;
      17'd57143: data = 8'h0a;
      17'd57144: data = 8'h05;
      17'd57145: data = 8'hd8;
      17'd57146: data = 8'h01;
      17'd57147: data = 8'he4;
      17'd57148: data = 8'hd8;
      17'd57149: data = 8'h04;
      17'd57150: data = 8'hdb;
      17'd57151: data = 8'hed;
      17'd57152: data = 8'hfe;
      17'd57153: data = 8'hd2;
      17'd57154: data = 8'hf4;
      17'd57155: data = 8'he4;
      17'd57156: data = 8'hcd;
      17'd57157: data = 8'hec;
      17'd57158: data = 8'hcd;
      17'd57159: data = 8'hc2;
      17'd57160: data = 8'hda;
      17'd57161: data = 8'hc2;
      17'd57162: data = 8'hd1;
      17'd57163: data = 8'he2;
      17'd57164: data = 8'hcd;
      17'd57165: data = 8'he5;
      17'd57166: data = 8'he4;
      17'd57167: data = 8'hdc;
      17'd57168: data = 8'hf5;
      17'd57169: data = 8'hec;
      17'd57170: data = 8'hed;
      17'd57171: data = 8'h04;
      17'd57172: data = 8'hf9;
      17'd57173: data = 8'h04;
      17'd57174: data = 8'h0a;
      17'd57175: data = 8'hfe;
      17'd57176: data = 8'h12;
      17'd57177: data = 8'h0c;
      17'd57178: data = 8'h0a;
      17'd57179: data = 8'h1e;
      17'd57180: data = 8'h12;
      17'd57181: data = 8'h15;
      17'd57182: data = 8'h29;
      17'd57183: data = 8'h22;
      17'd57184: data = 8'h26;
      17'd57185: data = 8'h2d;
      17'd57186: data = 8'h27;
      17'd57187: data = 8'h29;
      17'd57188: data = 8'h1b;
      17'd57189: data = 8'h1e;
      17'd57190: data = 8'h22;
      17'd57191: data = 8'h13;
      17'd57192: data = 8'h1a;
      17'd57193: data = 8'h1b;
      17'd57194: data = 8'h12;
      17'd57195: data = 8'h11;
      17'd57196: data = 8'h13;
      17'd57197: data = 8'h11;
      17'd57198: data = 8'h0d;
      17'd57199: data = 8'h0a;
      17'd57200: data = 8'h0c;
      17'd57201: data = 8'h05;
      17'd57202: data = 8'hfe;
      17'd57203: data = 8'h01;
      17'd57204: data = 8'hfd;
      17'd57205: data = 8'hfa;
      17'd57206: data = 8'hf5;
      17'd57207: data = 8'hf6;
      17'd57208: data = 8'hf4;
      17'd57209: data = 8'hf2;
      17'd57210: data = 8'hf2;
      17'd57211: data = 8'hf5;
      17'd57212: data = 8'hf9;
      17'd57213: data = 8'hfa;
      17'd57214: data = 8'h00;
      17'd57215: data = 8'h00;
      17'd57216: data = 8'h00;
      17'd57217: data = 8'h01;
      17'd57218: data = 8'h04;
      17'd57219: data = 8'h04;
      17'd57220: data = 8'h01;
      17'd57221: data = 8'h04;
      17'd57222: data = 8'h06;
      17'd57223: data = 8'h04;
      17'd57224: data = 8'h05;
      17'd57225: data = 8'h06;
      17'd57226: data = 8'h05;
      17'd57227: data = 8'h06;
      17'd57228: data = 8'h0a;
      17'd57229: data = 8'h0a;
      17'd57230: data = 8'h0a;
      17'd57231: data = 8'h09;
      17'd57232: data = 8'h05;
      17'd57233: data = 8'h02;
      17'd57234: data = 8'hfe;
      17'd57235: data = 8'hfe;
      17'd57236: data = 8'hfe;
      17'd57237: data = 8'hfd;
      17'd57238: data = 8'h01;
      17'd57239: data = 8'h04;
      17'd57240: data = 8'h02;
      17'd57241: data = 8'h04;
      17'd57242: data = 8'h01;
      17'd57243: data = 8'hfe;
      17'd57244: data = 8'hfa;
      17'd57245: data = 8'hf4;
      17'd57246: data = 8'hf2;
      17'd57247: data = 8'hf2;
      17'd57248: data = 8'hf2;
      17'd57249: data = 8'hf2;
      17'd57250: data = 8'hf2;
      17'd57251: data = 8'hf2;
      17'd57252: data = 8'hef;
      17'd57253: data = 8'heb;
      17'd57254: data = 8'he9;
      17'd57255: data = 8'he5;
      17'd57256: data = 8'he3;
      17'd57257: data = 8'he4;
      17'd57258: data = 8'he3;
      17'd57259: data = 8'he3;
      17'd57260: data = 8'he4;
      17'd57261: data = 8'he4;
      17'd57262: data = 8'he3;
      17'd57263: data = 8'he3;
      17'd57264: data = 8'he5;
      17'd57265: data = 8'he9;
      17'd57266: data = 8'he5;
      17'd57267: data = 8'he9;
      17'd57268: data = 8'hed;
      17'd57269: data = 8'hed;
      17'd57270: data = 8'hed;
      17'd57271: data = 8'hf1;
      17'd57272: data = 8'hf2;
      17'd57273: data = 8'hf1;
      17'd57274: data = 8'hed;
      17'd57275: data = 8'hf2;
      17'd57276: data = 8'hf1;
      17'd57277: data = 8'hf1;
      17'd57278: data = 8'hf5;
      17'd57279: data = 8'hf4;
      17'd57280: data = 8'hf4;
      17'd57281: data = 8'hf4;
      17'd57282: data = 8'hf4;
      17'd57283: data = 8'hf9;
      17'd57284: data = 8'hf9;
      17'd57285: data = 8'hfa;
      17'd57286: data = 8'h02;
      17'd57287: data = 8'h00;
      17'd57288: data = 8'hfd;
      17'd57289: data = 8'hfe;
      17'd57290: data = 8'hfd;
      17'd57291: data = 8'hfe;
      17'd57292: data = 8'h02;
      17'd57293: data = 8'h05;
      17'd57294: data = 8'h09;
      17'd57295: data = 8'h0c;
      17'd57296: data = 8'h0a;
      17'd57297: data = 8'h09;
      17'd57298: data = 8'h06;
      17'd57299: data = 8'h06;
      17'd57300: data = 8'h09;
      17'd57301: data = 8'h0a;
      17'd57302: data = 8'h09;
      17'd57303: data = 8'h0c;
      17'd57304: data = 8'h0c;
      17'd57305: data = 8'h09;
      17'd57306: data = 8'h0a;
      17'd57307: data = 8'h06;
      17'd57308: data = 8'h0a;
      17'd57309: data = 8'h0a;
      17'd57310: data = 8'h06;
      17'd57311: data = 8'h0a;
      17'd57312: data = 8'h09;
      17'd57313: data = 8'h09;
      17'd57314: data = 8'h0c;
      17'd57315: data = 8'h09;
      17'd57316: data = 8'h09;
      17'd57317: data = 8'h06;
      17'd57318: data = 8'h04;
      17'd57319: data = 8'h06;
      17'd57320: data = 8'h06;
      17'd57321: data = 8'h04;
      17'd57322: data = 8'h09;
      17'd57323: data = 8'h05;
      17'd57324: data = 8'h05;
      17'd57325: data = 8'h0a;
      17'd57326: data = 8'h06;
      17'd57327: data = 8'h05;
      17'd57328: data = 8'h04;
      17'd57329: data = 8'h02;
      17'd57330: data = 8'h09;
      17'd57331: data = 8'h04;
      17'd57332: data = 8'h02;
      17'd57333: data = 8'h05;
      17'd57334: data = 8'h09;
      17'd57335: data = 8'h0c;
      17'd57336: data = 8'h0c;
      17'd57337: data = 8'h06;
      17'd57338: data = 8'h00;
      17'd57339: data = 8'hfd;
      17'd57340: data = 8'hfd;
      17'd57341: data = 8'hfd;
      17'd57342: data = 8'hfe;
      17'd57343: data = 8'h05;
      17'd57344: data = 8'h09;
      17'd57345: data = 8'h05;
      17'd57346: data = 8'h0c;
      17'd57347: data = 8'h0a;
      17'd57348: data = 8'h01;
      17'd57349: data = 8'h00;
      17'd57350: data = 8'hfe;
      17'd57351: data = 8'h05;
      17'd57352: data = 8'h0d;
      17'd57353: data = 8'h0e;
      17'd57354: data = 8'h11;
      17'd57355: data = 8'h12;
      17'd57356: data = 8'h0d;
      17'd57357: data = 8'h0a;
      17'd57358: data = 8'h09;
      17'd57359: data = 8'h05;
      17'd57360: data = 8'h09;
      17'd57361: data = 8'h0c;
      17'd57362: data = 8'h0e;
      17'd57363: data = 8'h13;
      17'd57364: data = 8'h12;
      17'd57365: data = 8'h0e;
      17'd57366: data = 8'h0c;
      17'd57367: data = 8'h0a;
      17'd57368: data = 8'h09;
      17'd57369: data = 8'h05;
      17'd57370: data = 8'h04;
      17'd57371: data = 8'h06;
      17'd57372: data = 8'h05;
      17'd57373: data = 8'h05;
      17'd57374: data = 8'h04;
      17'd57375: data = 8'h04;
      17'd57376: data = 8'h01;
      17'd57377: data = 8'hfe;
      17'd57378: data = 8'h00;
      17'd57379: data = 8'h01;
      17'd57380: data = 8'h04;
      17'd57381: data = 8'h00;
      17'd57382: data = 8'hfc;
      17'd57383: data = 8'hfc;
      17'd57384: data = 8'hf5;
      17'd57385: data = 8'hf2;
      17'd57386: data = 8'hf1;
      17'd57387: data = 8'hef;
      17'd57388: data = 8'hf1;
      17'd57389: data = 8'hf2;
      17'd57390: data = 8'hf2;
      17'd57391: data = 8'hf1;
      17'd57392: data = 8'hef;
      17'd57393: data = 8'hec;
      17'd57394: data = 8'hed;
      17'd57395: data = 8'hec;
      17'd57396: data = 8'hef;
      17'd57397: data = 8'hf2;
      17'd57398: data = 8'hf5;
      17'd57399: data = 8'hf5;
      17'd57400: data = 8'hf5;
      17'd57401: data = 8'hf9;
      17'd57402: data = 8'hf6;
      17'd57403: data = 8'hf4;
      17'd57404: data = 8'hf4;
      17'd57405: data = 8'hf5;
      17'd57406: data = 8'hf4;
      17'd57407: data = 8'hf4;
      17'd57408: data = 8'hf6;
      17'd57409: data = 8'hf9;
      17'd57410: data = 8'hf9;
      17'd57411: data = 8'hf9;
      17'd57412: data = 8'hf9;
      17'd57413: data = 8'hf5;
      17'd57414: data = 8'hf6;
      17'd57415: data = 8'hf6;
      17'd57416: data = 8'hfa;
      17'd57417: data = 8'hfe;
      17'd57418: data = 8'h01;
      17'd57419: data = 8'hfe;
      17'd57420: data = 8'hfe;
      17'd57421: data = 8'hfe;
      17'd57422: data = 8'hfa;
      17'd57423: data = 8'hfe;
      17'd57424: data = 8'hfe;
      17'd57425: data = 8'h00;
      17'd57426: data = 8'h00;
      17'd57427: data = 8'h02;
      17'd57428: data = 8'h04;
      17'd57429: data = 8'h05;
      17'd57430: data = 8'h09;
      17'd57431: data = 8'h0a;
      17'd57432: data = 8'h09;
      17'd57433: data = 8'h0a;
      17'd57434: data = 8'h09;
      17'd57435: data = 8'h06;
      17'd57436: data = 8'h09;
      17'd57437: data = 8'h09;
      17'd57438: data = 8'h0a;
      17'd57439: data = 8'h0a;
      17'd57440: data = 8'h0c;
      17'd57441: data = 8'h0a;
      17'd57442: data = 8'h0a;
      17'd57443: data = 8'h09;
      17'd57444: data = 8'h09;
      17'd57445: data = 8'h0c;
      17'd57446: data = 8'h0c;
      17'd57447: data = 8'h0c;
      17'd57448: data = 8'h0c;
      17'd57449: data = 8'h0c;
      17'd57450: data = 8'h0d;
      17'd57451: data = 8'h0a;
      17'd57452: data = 8'h05;
      17'd57453: data = 8'h0a;
      17'd57454: data = 8'h04;
      17'd57455: data = 8'h02;
      17'd57456: data = 8'h02;
      17'd57457: data = 8'h00;
      17'd57458: data = 8'h02;
      17'd57459: data = 8'h04;
      17'd57460: data = 8'h04;
      17'd57461: data = 8'h04;
      17'd57462: data = 8'h01;
      17'd57463: data = 8'h02;
      17'd57464: data = 8'h01;
      17'd57465: data = 8'h01;
      17'd57466: data = 8'h02;
      17'd57467: data = 8'h04;
      17'd57468: data = 8'h02;
      17'd57469: data = 8'h04;
      17'd57470: data = 8'h04;
      17'd57471: data = 8'h01;
      17'd57472: data = 8'hfe;
      17'd57473: data = 8'h00;
      17'd57474: data = 8'h00;
      17'd57475: data = 8'h00;
      17'd57476: data = 8'h01;
      17'd57477: data = 8'hfe;
      17'd57478: data = 8'h01;
      17'd57479: data = 8'h01;
      17'd57480: data = 8'hfe;
      17'd57481: data = 8'h00;
      17'd57482: data = 8'h01;
      17'd57483: data = 8'hfe;
      17'd57484: data = 8'hfc;
      17'd57485: data = 8'hf9;
      17'd57486: data = 8'hf9;
      17'd57487: data = 8'hf5;
      17'd57488: data = 8'hf9;
      17'd57489: data = 8'hfc;
      17'd57490: data = 8'hf5;
      17'd57491: data = 8'hf4;
      17'd57492: data = 8'hf9;
      17'd57493: data = 8'hf5;
      17'd57494: data = 8'hf5;
      17'd57495: data = 8'hf5;
      17'd57496: data = 8'hf4;
      17'd57497: data = 8'hf4;
      17'd57498: data = 8'hef;
      17'd57499: data = 8'hec;
      17'd57500: data = 8'hec;
      17'd57501: data = 8'hec;
      17'd57502: data = 8'hed;
      17'd57503: data = 8'hef;
      17'd57504: data = 8'hef;
      17'd57505: data = 8'hec;
      17'd57506: data = 8'he9;
      17'd57507: data = 8'he7;
      17'd57508: data = 8'he7;
      17'd57509: data = 8'he9;
      17'd57510: data = 8'heb;
      17'd57511: data = 8'heb;
      17'd57512: data = 8'hed;
      17'd57513: data = 8'he7;
      17'd57514: data = 8'he9;
      17'd57515: data = 8'heb;
      17'd57516: data = 8'heb;
      17'd57517: data = 8'heb;
      17'd57518: data = 8'hed;
      17'd57519: data = 8'hf1;
      17'd57520: data = 8'hf1;
      17'd57521: data = 8'hf1;
      17'd57522: data = 8'hf1;
      17'd57523: data = 8'hef;
      17'd57524: data = 8'hf1;
      17'd57525: data = 8'hf4;
      17'd57526: data = 8'hf6;
      17'd57527: data = 8'hfa;
      17'd57528: data = 8'hfa;
      17'd57529: data = 8'hfa;
      17'd57530: data = 8'hfc;
      17'd57531: data = 8'hfd;
      17'd57532: data = 8'hfe;
      17'd57533: data = 8'hfe;
      17'd57534: data = 8'h01;
      17'd57535: data = 8'h04;
      17'd57536: data = 8'h05;
      17'd57537: data = 8'h0a;
      17'd57538: data = 8'h0a;
      17'd57539: data = 8'h0c;
      17'd57540: data = 8'h0c;
      17'd57541: data = 8'h09;
      17'd57542: data = 8'h0a;
      17'd57543: data = 8'h09;
      17'd57544: data = 8'h09;
      17'd57545: data = 8'h0c;
      17'd57546: data = 8'h0e;
      17'd57547: data = 8'h12;
      17'd57548: data = 8'h13;
      17'd57549: data = 8'h12;
      17'd57550: data = 8'h0d;
      17'd57551: data = 8'h0a;
      17'd57552: data = 8'h0a;
      17'd57553: data = 8'h0e;
      17'd57554: data = 8'h0d;
      17'd57555: data = 8'h0d;
      17'd57556: data = 8'h12;
      17'd57557: data = 8'h15;
      17'd57558: data = 8'h13;
      17'd57559: data = 8'h11;
      17'd57560: data = 8'h11;
      17'd57561: data = 8'h12;
      17'd57562: data = 8'h0d;
      17'd57563: data = 8'h0a;
      17'd57564: data = 8'h0c;
      17'd57565: data = 8'h0e;
      17'd57566: data = 8'h0c;
      17'd57567: data = 8'h09;
      17'd57568: data = 8'h06;
      17'd57569: data = 8'h09;
      17'd57570: data = 8'h0c;
      17'd57571: data = 8'h05;
      17'd57572: data = 8'h06;
      17'd57573: data = 8'h0a;
      17'd57574: data = 8'h05;
      17'd57575: data = 8'h04;
      17'd57576: data = 8'h09;
      17'd57577: data = 8'h05;
      17'd57578: data = 8'h01;
      17'd57579: data = 8'h06;
      17'd57580: data = 8'h12;
      17'd57581: data = 8'h11;
      17'd57582: data = 8'h0c;
      17'd57583: data = 8'h0a;
      17'd57584: data = 8'h0c;
      17'd57585: data = 8'h0a;
      17'd57586: data = 8'h02;
      17'd57587: data = 8'h04;
      17'd57588: data = 8'h0c;
      17'd57589: data = 8'h0d;
      17'd57590: data = 8'h04;
      17'd57591: data = 8'h02;
      17'd57592: data = 8'h09;
      17'd57593: data = 8'h01;
      17'd57594: data = 8'hfc;
      17'd57595: data = 8'hfe;
      17'd57596: data = 8'h00;
      17'd57597: data = 8'h00;
      17'd57598: data = 8'h00;
      17'd57599: data = 8'h01;
      17'd57600: data = 8'h01;
      17'd57601: data = 8'h00;
      17'd57602: data = 8'hfd;
      17'd57603: data = 8'hfd;
      17'd57604: data = 8'h00;
      17'd57605: data = 8'hfc;
      17'd57606: data = 8'hf6;
      17'd57607: data = 8'hfc;
      17'd57608: data = 8'hfc;
      17'd57609: data = 8'hf6;
      17'd57610: data = 8'hf6;
      17'd57611: data = 8'hf5;
      17'd57612: data = 8'hf2;
      17'd57613: data = 8'hf2;
      17'd57614: data = 8'hf1;
      17'd57615: data = 8'hf1;
      17'd57616: data = 8'hf1;
      17'd57617: data = 8'hf1;
      17'd57618: data = 8'hef;
      17'd57619: data = 8'hed;
      17'd57620: data = 8'hed;
      17'd57621: data = 8'hef;
      17'd57622: data = 8'heb;
      17'd57623: data = 8'hec;
      17'd57624: data = 8'he9;
      17'd57625: data = 8'heb;
      17'd57626: data = 8'hf2;
      17'd57627: data = 8'hf1;
      17'd57628: data = 8'hef;
      17'd57629: data = 8'hf1;
      17'd57630: data = 8'hf1;
      17'd57631: data = 8'hef;
      17'd57632: data = 8'hf4;
      17'd57633: data = 8'hf4;
      17'd57634: data = 8'hf6;
      17'd57635: data = 8'hfa;
      17'd57636: data = 8'hf6;
      17'd57637: data = 8'hf6;
      17'd57638: data = 8'hf5;
      17'd57639: data = 8'hf2;
      17'd57640: data = 8'hf5;
      17'd57641: data = 8'hfc;
      17'd57642: data = 8'hfe;
      17'd57643: data = 8'h00;
      17'd57644: data = 8'h01;
      17'd57645: data = 8'h09;
      17'd57646: data = 8'h05;
      17'd57647: data = 8'h04;
      17'd57648: data = 8'h0c;
      17'd57649: data = 8'h0d;
      17'd57650: data = 8'h0d;
      17'd57651: data = 8'h0e;
      17'd57652: data = 8'h11;
      17'd57653: data = 8'h12;
      17'd57654: data = 8'h0e;
      17'd57655: data = 8'h0e;
      17'd57656: data = 8'h11;
      17'd57657: data = 8'h12;
      17'd57658: data = 8'h0e;
      17'd57659: data = 8'h0d;
      17'd57660: data = 8'h0e;
      17'd57661: data = 8'h0d;
      17'd57662: data = 8'h0d;
      17'd57663: data = 8'h0a;
      17'd57664: data = 8'h0e;
      17'd57665: data = 8'h11;
      17'd57666: data = 8'h0a;
      17'd57667: data = 8'h0c;
      17'd57668: data = 8'h0d;
      17'd57669: data = 8'h0d;
      17'd57670: data = 8'h0e;
      17'd57671: data = 8'h0d;
      17'd57672: data = 8'h0c;
      17'd57673: data = 8'h0c;
      17'd57674: data = 8'h09;
      17'd57675: data = 8'h05;
      17'd57676: data = 8'h04;
      17'd57677: data = 8'h05;
      17'd57678: data = 8'h06;
      17'd57679: data = 8'h06;
      17'd57680: data = 8'h04;
      17'd57681: data = 8'h05;
      17'd57682: data = 8'h05;
      17'd57683: data = 8'h02;
      17'd57684: data = 8'h05;
      17'd57685: data = 8'h06;
      17'd57686: data = 8'h05;
      17'd57687: data = 8'h04;
      17'd57688: data = 8'h02;
      17'd57689: data = 8'h04;
      17'd57690: data = 8'h05;
      17'd57691: data = 8'h01;
      17'd57692: data = 8'hfe;
      17'd57693: data = 8'h01;
      17'd57694: data = 8'h04;
      17'd57695: data = 8'h04;
      17'd57696: data = 8'h00;
      17'd57697: data = 8'hfd;
      17'd57698: data = 8'h02;
      17'd57699: data = 8'h02;
      17'd57700: data = 8'h01;
      17'd57701: data = 8'h00;
      17'd57702: data = 8'hfe;
      17'd57703: data = 8'hfe;
      17'd57704: data = 8'hfa;
      17'd57705: data = 8'hf6;
      17'd57706: data = 8'hf9;
      17'd57707: data = 8'hf4;
      17'd57708: data = 8'hf4;
      17'd57709: data = 8'hf6;
      17'd57710: data = 8'hf2;
      17'd57711: data = 8'hf5;
      17'd57712: data = 8'hf1;
      17'd57713: data = 8'heb;
      17'd57714: data = 8'hed;
      17'd57715: data = 8'hec;
      17'd57716: data = 8'he9;
      17'd57717: data = 8'hec;
      17'd57718: data = 8'hef;
      17'd57719: data = 8'hef;
      17'd57720: data = 8'hec;
      17'd57721: data = 8'heb;
      17'd57722: data = 8'hed;
      17'd57723: data = 8'heb;
      17'd57724: data = 8'he7;
      17'd57725: data = 8'heb;
      17'd57726: data = 8'heb;
      17'd57727: data = 8'he9;
      17'd57728: data = 8'heb;
      17'd57729: data = 8'he7;
      17'd57730: data = 8'he9;
      17'd57731: data = 8'he7;
      17'd57732: data = 8'he3;
      17'd57733: data = 8'he3;
      17'd57734: data = 8'he7;
      17'd57735: data = 8'he9;
      17'd57736: data = 8'he9;
      17'd57737: data = 8'he9;
      17'd57738: data = 8'he9;
      17'd57739: data = 8'hed;
      17'd57740: data = 8'hec;
      17'd57741: data = 8'heb;
      17'd57742: data = 8'hec;
      17'd57743: data = 8'hef;
      17'd57744: data = 8'hef;
      17'd57745: data = 8'hf1;
      17'd57746: data = 8'hf2;
      17'd57747: data = 8'hf4;
      17'd57748: data = 8'hf4;
      17'd57749: data = 8'hf5;
      17'd57750: data = 8'hf9;
      17'd57751: data = 8'hf9;
      17'd57752: data = 8'hfc;
      17'd57753: data = 8'hfe;
      17'd57754: data = 8'hfd;
      17'd57755: data = 8'h00;
      17'd57756: data = 8'h02;
      17'd57757: data = 8'h01;
      17'd57758: data = 8'h01;
      17'd57759: data = 8'h05;
      17'd57760: data = 8'h05;
      17'd57761: data = 8'h04;
      17'd57762: data = 8'h09;
      17'd57763: data = 8'h0a;
      17'd57764: data = 8'h0a;
      17'd57765: data = 8'h0a;
      17'd57766: data = 8'h09;
      17'd57767: data = 8'h0e;
      17'd57768: data = 8'h0e;
      17'd57769: data = 8'h09;
      17'd57770: data = 8'h0c;
      17'd57771: data = 8'h12;
      17'd57772: data = 8'h16;
      17'd57773: data = 8'h0e;
      17'd57774: data = 8'h06;
      17'd57775: data = 8'h0d;
      17'd57776: data = 8'h0d;
      17'd57777: data = 8'h0c;
      17'd57778: data = 8'h0a;
      17'd57779: data = 8'h09;
      17'd57780: data = 8'h12;
      17'd57781: data = 8'h1c;
      17'd57782: data = 8'h19;
      17'd57783: data = 8'h13;
      17'd57784: data = 8'h16;
      17'd57785: data = 8'h11;
      17'd57786: data = 8'h12;
      17'd57787: data = 8'h0d;
      17'd57788: data = 8'h02;
      17'd57789: data = 8'h04;
      17'd57790: data = 8'h0e;
      17'd57791: data = 8'h0d;
      17'd57792: data = 8'h05;
      17'd57793: data = 8'h05;
      17'd57794: data = 8'h06;
      17'd57795: data = 8'h0c;
      17'd57796: data = 8'h06;
      17'd57797: data = 8'h05;
      17'd57798: data = 8'h05;
      17'd57799: data = 8'h0c;
      17'd57800: data = 8'h11;
      17'd57801: data = 8'h06;
      17'd57802: data = 8'h06;
      17'd57803: data = 8'h0e;
      17'd57804: data = 8'h0d;
      17'd57805: data = 8'h0e;
      17'd57806: data = 8'h0e;
      17'd57807: data = 8'h06;
      17'd57808: data = 8'h06;
      17'd57809: data = 8'h0a;
      17'd57810: data = 8'h05;
      17'd57811: data = 8'h05;
      17'd57812: data = 8'h06;
      17'd57813: data = 8'h05;
      17'd57814: data = 8'h09;
      17'd57815: data = 8'h05;
      17'd57816: data = 8'h02;
      17'd57817: data = 8'h02;
      17'd57818: data = 8'h01;
      17'd57819: data = 8'h02;
      17'd57820: data = 8'hfe;
      17'd57821: data = 8'hfe;
      17'd57822: data = 8'h01;
      17'd57823: data = 8'hfe;
      17'd57824: data = 8'h01;
      17'd57825: data = 8'hfe;
      17'd57826: data = 8'h00;
      17'd57827: data = 8'h01;
      17'd57828: data = 8'h01;
      17'd57829: data = 8'hfd;
      17'd57830: data = 8'hfc;
      17'd57831: data = 8'hfc;
      17'd57832: data = 8'hfc;
      17'd57833: data = 8'hfd;
      17'd57834: data = 8'hf5;
      17'd57835: data = 8'hf2;
      17'd57836: data = 8'hf2;
      17'd57837: data = 8'hef;
      17'd57838: data = 8'hec;
      17'd57839: data = 8'heb;
      17'd57840: data = 8'hec;
      17'd57841: data = 8'hed;
      17'd57842: data = 8'hec;
      17'd57843: data = 8'he9;
      17'd57844: data = 8'hec;
      17'd57845: data = 8'heb;
      17'd57846: data = 8'hed;
      17'd57847: data = 8'hf1;
      17'd57848: data = 8'hef;
      17'd57849: data = 8'hef;
      17'd57850: data = 8'hed;
      17'd57851: data = 8'hef;
      17'd57852: data = 8'hf4;
      17'd57853: data = 8'hf1;
      17'd57854: data = 8'hf1;
      17'd57855: data = 8'hf5;
      17'd57856: data = 8'hf2;
      17'd57857: data = 8'hf6;
      17'd57858: data = 8'hf6;
      17'd57859: data = 8'hf4;
      17'd57860: data = 8'hfd;
      17'd57861: data = 8'hfe;
      17'd57862: data = 8'h00;
      17'd57863: data = 8'h02;
      17'd57864: data = 8'h00;
      17'd57865: data = 8'h02;
      17'd57866: data = 8'h05;
      17'd57867: data = 8'h05;
      17'd57868: data = 8'h0c;
      17'd57869: data = 8'h11;
      17'd57870: data = 8'h11;
      17'd57871: data = 8'h12;
      17'd57872: data = 8'h12;
      17'd57873: data = 8'h13;
      17'd57874: data = 8'h15;
      17'd57875: data = 8'h16;
      17'd57876: data = 8'h19;
      17'd57877: data = 8'h15;
      17'd57878: data = 8'h12;
      17'd57879: data = 8'h15;
      17'd57880: data = 8'h13;
      17'd57881: data = 8'h11;
      17'd57882: data = 8'h11;
      17'd57883: data = 8'h11;
      17'd57884: data = 8'h0e;
      17'd57885: data = 8'h11;
      17'd57886: data = 8'h0e;
      17'd57887: data = 8'h0c;
      17'd57888: data = 8'h0e;
      17'd57889: data = 8'h0e;
      17'd57890: data = 8'h0d;
      17'd57891: data = 8'h0c;
      17'd57892: data = 8'h0a;
      17'd57893: data = 8'h09;
      17'd57894: data = 8'h06;
      17'd57895: data = 8'h05;
      17'd57896: data = 8'h05;
      17'd57897: data = 8'h05;
      17'd57898: data = 8'h06;
      17'd57899: data = 8'h06;
      17'd57900: data = 8'h05;
      17'd57901: data = 8'h02;
      17'd57902: data = 8'h04;
      17'd57903: data = 8'h04;
      17'd57904: data = 8'h04;
      17'd57905: data = 8'h02;
      17'd57906: data = 8'h01;
      17'd57907: data = 8'h00;
      17'd57908: data = 8'h00;
      17'd57909: data = 8'h01;
      17'd57910: data = 8'h02;
      17'd57911: data = 8'h04;
      17'd57912: data = 8'h04;
      17'd57913: data = 8'h04;
      17'd57914: data = 8'h01;
      17'd57915: data = 8'h02;
      17'd57916: data = 8'h01;
      17'd57917: data = 8'hfe;
      17'd57918: data = 8'h01;
      17'd57919: data = 8'h06;
      17'd57920: data = 8'h06;
      17'd57921: data = 8'h02;
      17'd57922: data = 8'h01;
      17'd57923: data = 8'h02;
      17'd57924: data = 8'hfd;
      17'd57925: data = 8'hfa;
      17'd57926: data = 8'hfa;
      17'd57927: data = 8'hf9;
      17'd57928: data = 8'hf9;
      17'd57929: data = 8'hfa;
      17'd57930: data = 8'hf9;
      17'd57931: data = 8'hfa;
      17'd57932: data = 8'hfa;
      17'd57933: data = 8'hf4;
      17'd57934: data = 8'hf2;
      17'd57935: data = 8'hef;
      17'd57936: data = 8'hed;
      17'd57937: data = 8'hec;
      17'd57938: data = 8'hec;
      17'd57939: data = 8'hec;
      17'd57940: data = 8'hed;
      17'd57941: data = 8'he9;
      17'd57942: data = 8'he9;
      17'd57943: data = 8'he9;
      17'd57944: data = 8'he5;
      17'd57945: data = 8'he7;
      17'd57946: data = 8'he7;
      17'd57947: data = 8'he7;
      17'd57948: data = 8'he7;
      17'd57949: data = 8'he7;
      17'd57950: data = 8'he5;
      17'd57951: data = 8'he3;
      17'd57952: data = 8'he0;
      17'd57953: data = 8'he2;
      17'd57954: data = 8'he0;
      17'd57955: data = 8'he2;
      17'd57956: data = 8'he3;
      17'd57957: data = 8'he0;
      17'd57958: data = 8'hde;
      17'd57959: data = 8'he0;
      17'd57960: data = 8'he0;
      17'd57961: data = 8'he3;
      17'd57962: data = 8'he9;
      17'd57963: data = 8'he9;
      17'd57964: data = 8'he7;
      17'd57965: data = 8'he7;
      17'd57966: data = 8'heb;
      17'd57967: data = 8'hef;
      17'd57968: data = 8'hed;
      17'd57969: data = 8'hef;
      17'd57970: data = 8'hf2;
      17'd57971: data = 8'hf5;
      17'd57972: data = 8'hf6;
      17'd57973: data = 8'hf6;
      17'd57974: data = 8'hfa;
      17'd57975: data = 8'hfc;
      17'd57976: data = 8'hfd;
      17'd57977: data = 8'h01;
      17'd57978: data = 8'h02;
      17'd57979: data = 8'h02;
      17'd57980: data = 8'h04;
      17'd57981: data = 8'h04;
      17'd57982: data = 8'h06;
      17'd57983: data = 8'h0c;
      17'd57984: data = 8'h0d;
      17'd57985: data = 8'h0e;
      17'd57986: data = 8'h0d;
      17'd57987: data = 8'h09;
      17'd57988: data = 8'h0c;
      17'd57989: data = 8'h0e;
      17'd57990: data = 8'h0d;
      17'd57991: data = 8'h0c;
      17'd57992: data = 8'h12;
      17'd57993: data = 8'h13;
      17'd57994: data = 8'h15;
      17'd57995: data = 8'h15;
      17'd57996: data = 8'h15;
      17'd57997: data = 8'h13;
      17'd57998: data = 8'h12;
      17'd57999: data = 8'h12;
      17'd58000: data = 8'h11;
      17'd58001: data = 8'h0e;
      17'd58002: data = 8'h11;
      17'd58003: data = 8'h16;
      17'd58004: data = 8'h16;
      17'd58005: data = 8'h15;
      17'd58006: data = 8'h16;
      17'd58007: data = 8'h16;
      17'd58008: data = 8'h0e;
      17'd58009: data = 8'h0a;
      17'd58010: data = 8'h06;
      17'd58011: data = 8'h05;
      17'd58012: data = 8'h06;
      17'd58013: data = 8'h0a;
      17'd58014: data = 8'h0e;
      17'd58015: data = 8'h0a;
      17'd58016: data = 8'h09;
      17'd58017: data = 8'h06;
      17'd58018: data = 8'h05;
      17'd58019: data = 8'h01;
      17'd58020: data = 8'h04;
      17'd58021: data = 8'h0a;
      17'd58022: data = 8'h0d;
      17'd58023: data = 8'h0d;
      17'd58024: data = 8'h0d;
      17'd58025: data = 8'h0e;
      17'd58026: data = 8'h0e;
      17'd58027: data = 8'h0a;
      17'd58028: data = 8'h0a;
      17'd58029: data = 8'h0c;
      17'd58030: data = 8'h0a;
      17'd58031: data = 8'h0a;
      17'd58032: data = 8'h0c;
      17'd58033: data = 8'h09;
      17'd58034: data = 8'h05;
      17'd58035: data = 8'h06;
      17'd58036: data = 8'h09;
      17'd58037: data = 8'h06;
      17'd58038: data = 8'h05;
      17'd58039: data = 8'h05;
      17'd58040: data = 8'h09;
      17'd58041: data = 8'h06;
      17'd58042: data = 8'h04;
      17'd58043: data = 8'h02;
      17'd58044: data = 8'h04;
      17'd58045: data = 8'h02;
      17'd58046: data = 8'h00;
      17'd58047: data = 8'h01;
      17'd58048: data = 8'h04;
      17'd58049: data = 8'h02;
      17'd58050: data = 8'h02;
      17'd58051: data = 8'h01;
      17'd58052: data = 8'hfd;
      17'd58053: data = 8'hfc;
      17'd58054: data = 8'hfa;
      17'd58055: data = 8'hf9;
      17'd58056: data = 8'hf5;
      17'd58057: data = 8'hf1;
      17'd58058: data = 8'hf2;
      17'd58059: data = 8'hf1;
      17'd58060: data = 8'hec;
      17'd58061: data = 8'heb;
      17'd58062: data = 8'heb;
      17'd58063: data = 8'heb;
      17'd58064: data = 8'he7;
      17'd58065: data = 8'he7;
      17'd58066: data = 8'he9;
      17'd58067: data = 8'he9;
      17'd58068: data = 8'he5;
      17'd58069: data = 8'heb;
      17'd58070: data = 8'hec;
      17'd58071: data = 8'heb;
      17'd58072: data = 8'hec;
      17'd58073: data = 8'hec;
      17'd58074: data = 8'heb;
      17'd58075: data = 8'heb;
      17'd58076: data = 8'hec;
      17'd58077: data = 8'hed;
      17'd58078: data = 8'hf1;
      17'd58079: data = 8'hf1;
      17'd58080: data = 8'hf1;
      17'd58081: data = 8'hf4;
      17'd58082: data = 8'hf2;
      17'd58083: data = 8'hf2;
      17'd58084: data = 8'hfc;
      17'd58085: data = 8'hfe;
      17'd58086: data = 8'hfd;
      17'd58087: data = 8'h00;
      17'd58088: data = 8'h04;
      17'd58089: data = 8'h06;
      17'd58090: data = 8'h05;
      17'd58091: data = 8'h09;
      17'd58092: data = 8'h0c;
      17'd58093: data = 8'h0e;
      17'd58094: data = 8'h0e;
      17'd58095: data = 8'h11;
      17'd58096: data = 8'h13;
      17'd58097: data = 8'h13;
      17'd58098: data = 8'h13;
      17'd58099: data = 8'h12;
      17'd58100: data = 8'h15;
      17'd58101: data = 8'h15;
      17'd58102: data = 8'h11;
      17'd58103: data = 8'h15;
      17'd58104: data = 8'h15;
      17'd58105: data = 8'h13;
      17'd58106: data = 8'h13;
      17'd58107: data = 8'h12;
      17'd58108: data = 8'h13;
      17'd58109: data = 8'h11;
      17'd58110: data = 8'h0d;
      17'd58111: data = 8'h11;
      17'd58112: data = 8'h11;
      17'd58113: data = 8'h11;
      17'd58114: data = 8'h0e;
      17'd58115: data = 8'h11;
      17'd58116: data = 8'h0e;
      17'd58117: data = 8'h0a;
      17'd58118: data = 8'h0a;
      17'd58119: data = 8'h09;
      17'd58120: data = 8'h04;
      17'd58121: data = 8'h04;
      17'd58122: data = 8'h05;
      17'd58123: data = 8'h04;
      17'd58124: data = 8'h05;
      17'd58125: data = 8'h05;
      17'd58126: data = 8'h05;
      17'd58127: data = 8'h01;
      17'd58128: data = 8'h00;
      17'd58129: data = 8'hfd;
      17'd58130: data = 8'hfe;
      17'd58131: data = 8'h01;
      17'd58132: data = 8'h00;
      17'd58133: data = 8'hfe;
      17'd58134: data = 8'h01;
      17'd58135: data = 8'h01;
      17'd58136: data = 8'hfe;
      17'd58137: data = 8'hfd;
      17'd58138: data = 8'hfe;
      17'd58139: data = 8'hfd;
      17'd58140: data = 8'hfd;
      17'd58141: data = 8'h01;
      17'd58142: data = 8'h02;
      17'd58143: data = 8'h01;
      17'd58144: data = 8'h00;
      17'd58145: data = 8'hfd;
      17'd58146: data = 8'hfa;
      17'd58147: data = 8'hf6;
      17'd58148: data = 8'hf2;
      17'd58149: data = 8'hf5;
      17'd58150: data = 8'hf5;
      17'd58151: data = 8'hf6;
      17'd58152: data = 8'hf9;
      17'd58153: data = 8'hf4;
      17'd58154: data = 8'hf2;
      17'd58155: data = 8'hf1;
      17'd58156: data = 8'hf1;
      17'd58157: data = 8'hf2;
      17'd58158: data = 8'hf2;
      17'd58159: data = 8'hf2;
      17'd58160: data = 8'hf2;
      17'd58161: data = 8'hf2;
      17'd58162: data = 8'hef;
      17'd58163: data = 8'hed;
      17'd58164: data = 8'hec;
      17'd58165: data = 8'heb;
      17'd58166: data = 8'he9;
      17'd58167: data = 8'he9;
      17'd58168: data = 8'he9;
      17'd58169: data = 8'he9;
      17'd58170: data = 8'he7;
      17'd58171: data = 8'he9;
      17'd58172: data = 8'heb;
      17'd58173: data = 8'he9;
      17'd58174: data = 8'he5;
      17'd58175: data = 8'he2;
      17'd58176: data = 8'he0;
      17'd58177: data = 8'he0;
      17'd58178: data = 8'he0;
      17'd58179: data = 8'hde;
      17'd58180: data = 8'he0;
      17'd58181: data = 8'he0;
      17'd58182: data = 8'he0;
      17'd58183: data = 8'he0;
      17'd58184: data = 8'hde;
      17'd58185: data = 8'he2;
      17'd58186: data = 8'he7;
      17'd58187: data = 8'hed;
      17'd58188: data = 8'hec;
      17'd58189: data = 8'hed;
      17'd58190: data = 8'hec;
      17'd58191: data = 8'hec;
      17'd58192: data = 8'hef;
      17'd58193: data = 8'heb;
      17'd58194: data = 8'hed;
      17'd58195: data = 8'hed;
      17'd58196: data = 8'hf6;
      17'd58197: data = 8'hf6;
      17'd58198: data = 8'hf6;
      17'd58199: data = 8'hfd;
      17'd58200: data = 8'hfd;
      17'd58201: data = 8'h09;
      17'd58202: data = 8'h00;
      17'd58203: data = 8'h02;
      17'd58204: data = 8'hfd;
      17'd58205: data = 8'h05;
      17'd58206: data = 8'h0a;
      17'd58207: data = 8'h15;
      17'd58208: data = 8'h12;
      17'd58209: data = 8'h0c;
      17'd58210: data = 8'h0c;
      17'd58211: data = 8'h04;
      17'd58212: data = 8'h0d;
      17'd58213: data = 8'h05;
      17'd58214: data = 8'h15;
      17'd58215: data = 8'h19;
      17'd58216: data = 8'h27;
      17'd58217: data = 8'h1a;
      17'd58218: data = 8'h1c;
      17'd58219: data = 8'h0c;
      17'd58220: data = 8'h12;
      17'd58221: data = 8'h15;
      17'd58222: data = 8'h12;
      17'd58223: data = 8'h1f;
      17'd58224: data = 8'h19;
      17'd58225: data = 8'h1c;
      17'd58226: data = 8'h04;
      17'd58227: data = 8'hfe;
      17'd58228: data = 8'hfc;
      17'd58229: data = 8'h13;
      17'd58230: data = 8'h16;
      17'd58231: data = 8'h1a;
      17'd58232: data = 8'h04;
      17'd58233: data = 8'h04;
      17'd58234: data = 8'h05;
      17'd58235: data = 8'h06;
      17'd58236: data = 8'h12;
      17'd58237: data = 8'h13;
      17'd58238: data = 8'h16;
      17'd58239: data = 8'h02;
      17'd58240: data = 8'hfd;
      17'd58241: data = 8'hf2;
      17'd58242: data = 8'h04;
      17'd58243: data = 8'h0c;
      17'd58244: data = 8'h23;
      17'd58245: data = 8'h2d;
      17'd58246: data = 8'h22;
      17'd58247: data = 8'h0e;
      17'd58248: data = 8'h06;
      17'd58249: data = 8'h0c;
      17'd58250: data = 8'h0d;
      17'd58251: data = 8'h1b;
      17'd58252: data = 8'h19;
      17'd58253: data = 8'h23;
      17'd58254: data = 8'h0e;
      17'd58255: data = 8'h02;
      17'd58256: data = 8'hfd;
      17'd58257: data = 8'h06;
      17'd58258: data = 8'h0c;
      17'd58259: data = 8'h16;
      17'd58260: data = 8'h1c;
      17'd58261: data = 8'h09;
      17'd58262: data = 8'h02;
      17'd58263: data = 8'hfd;
      17'd58264: data = 8'h04;
      17'd58265: data = 8'h05;
      17'd58266: data = 8'h0d;
      17'd58267: data = 8'h05;
      17'd58268: data = 8'hfe;
      17'd58269: data = 8'he7;
      17'd58270: data = 8'he9;
      17'd58271: data = 8'hf6;
      17'd58272: data = 8'h02;
      17'd58273: data = 8'h09;
      17'd58274: data = 8'hfc;
      17'd58275: data = 8'hf4;
      17'd58276: data = 8'he2;
      17'd58277: data = 8'hdb;
      17'd58278: data = 8'he0;
      17'd58279: data = 8'hf2;
      17'd58280: data = 8'hf5;
      17'd58281: data = 8'hf1;
      17'd58282: data = 8'hed;
      17'd58283: data = 8'hd6;
      17'd58284: data = 8'hd6;
      17'd58285: data = 8'hd6;
      17'd58286: data = 8'he5;
      17'd58287: data = 8'hf4;
      17'd58288: data = 8'hf1;
      17'd58289: data = 8'hec;
      17'd58290: data = 8'hed;
      17'd58291: data = 8'he5;
      17'd58292: data = 8'he2;
      17'd58293: data = 8'hed;
      17'd58294: data = 8'hf1;
      17'd58295: data = 8'hf9;
      17'd58296: data = 8'hed;
      17'd58297: data = 8'hf2;
      17'd58298: data = 8'hf2;
      17'd58299: data = 8'hf6;
      17'd58300: data = 8'h01;
      17'd58301: data = 8'h0c;
      17'd58302: data = 8'h0c;
      17'd58303: data = 8'hfa;
      17'd58304: data = 8'hf6;
      17'd58305: data = 8'hf6;
      17'd58306: data = 8'h01;
      17'd58307: data = 8'h00;
      17'd58308: data = 8'h11;
      17'd58309: data = 8'h12;
      17'd58310: data = 8'h0c;
      17'd58311: data = 8'h04;
      17'd58312: data = 8'h01;
      17'd58313: data = 8'h0c;
      17'd58314: data = 8'h12;
      17'd58315: data = 8'h19;
      17'd58316: data = 8'h1b;
      17'd58317: data = 8'h19;
      17'd58318: data = 8'h0d;
      17'd58319: data = 8'h0c;
      17'd58320: data = 8'h0a;
      17'd58321: data = 8'h0a;
      17'd58322: data = 8'h0a;
      17'd58323: data = 8'h05;
      17'd58324: data = 8'h06;
      17'd58325: data = 8'h06;
      17'd58326: data = 8'h06;
      17'd58327: data = 8'h12;
      17'd58328: data = 8'h16;
      17'd58329: data = 8'h16;
      17'd58330: data = 8'h15;
      17'd58331: data = 8'h0d;
      17'd58332: data = 8'h06;
      17'd58333: data = 8'h05;
      17'd58334: data = 8'h09;
      17'd58335: data = 8'h0e;
      17'd58336: data = 8'h0d;
      17'd58337: data = 8'h06;
      17'd58338: data = 8'h09;
      17'd58339: data = 8'h04;
      17'd58340: data = 8'h04;
      17'd58341: data = 8'h06;
      17'd58342: data = 8'h0e;
      17'd58343: data = 8'h12;
      17'd58344: data = 8'h0d;
      17'd58345: data = 8'h0c;
      17'd58346: data = 8'h11;
      17'd58347: data = 8'h0e;
      17'd58348: data = 8'h06;
      17'd58349: data = 8'h05;
      17'd58350: data = 8'h01;
      17'd58351: data = 8'h01;
      17'd58352: data = 8'h04;
      17'd58353: data = 8'h02;
      17'd58354: data = 8'h09;
      17'd58355: data = 8'h0c;
      17'd58356: data = 8'h0c;
      17'd58357: data = 8'h0c;
      17'd58358: data = 8'h05;
      17'd58359: data = 8'h01;
      17'd58360: data = 8'h00;
      17'd58361: data = 8'h01;
      17'd58362: data = 8'h01;
      17'd58363: data = 8'h04;
      17'd58364: data = 8'h02;
      17'd58365: data = 8'hfe;
      17'd58366: data = 8'hfa;
      17'd58367: data = 8'hf4;
      17'd58368: data = 8'hf4;
      17'd58369: data = 8'hf4;
      17'd58370: data = 8'hf4;
      17'd58371: data = 8'hf6;
      17'd58372: data = 8'hf5;
      17'd58373: data = 8'hef;
      17'd58374: data = 8'hed;
      17'd58375: data = 8'heb;
      17'd58376: data = 8'hec;
      17'd58377: data = 8'he9;
      17'd58378: data = 8'he5;
      17'd58379: data = 8'he5;
      17'd58380: data = 8'he5;
      17'd58381: data = 8'he9;
      17'd58382: data = 8'he7;
      17'd58383: data = 8'he4;
      17'd58384: data = 8'he0;
      17'd58385: data = 8'hdc;
      17'd58386: data = 8'hdb;
      17'd58387: data = 8'hdc;
      17'd58388: data = 8'he3;
      17'd58389: data = 8'he4;
      17'd58390: data = 8'he5;
      17'd58391: data = 8'he4;
      17'd58392: data = 8'he4;
      17'd58393: data = 8'he7;
      17'd58394: data = 8'he3;
      17'd58395: data = 8'he3;
      17'd58396: data = 8'he2;
      17'd58397: data = 8'he0;
      17'd58398: data = 8'hde;
      17'd58399: data = 8'hde;
      17'd58400: data = 8'he3;
      17'd58401: data = 8'he4;
      17'd58402: data = 8'he9;
      17'd58403: data = 8'he9;
      17'd58404: data = 8'hec;
      17'd58405: data = 8'hed;
      17'd58406: data = 8'hf1;
      17'd58407: data = 8'hf4;
      17'd58408: data = 8'hf5;
      17'd58409: data = 8'hfc;
      17'd58410: data = 8'hf6;
      17'd58411: data = 8'hf5;
      17'd58412: data = 8'hf2;
      17'd58413: data = 8'hf5;
      17'd58414: data = 8'hf5;
      17'd58415: data = 8'hfe;
      17'd58416: data = 8'h06;
      17'd58417: data = 8'h09;
      17'd58418: data = 8'h0c;
      17'd58419: data = 8'h09;
      17'd58420: data = 8'h0c;
      17'd58421: data = 8'h01;
      17'd58422: data = 8'h05;
      17'd58423: data = 8'h09;
      17'd58424: data = 8'h11;
      17'd58425: data = 8'h11;
      17'd58426: data = 8'h0a;
      17'd58427: data = 8'h1a;
      17'd58428: data = 8'h06;
      17'd58429: data = 8'h04;
      17'd58430: data = 8'h16;
      17'd58431: data = 8'h13;
      17'd58432: data = 8'hfd;
      17'd58433: data = 8'h0c;
      17'd58434: data = 8'h0e;
      17'd58435: data = 8'h0c;
      17'd58436: data = 8'h16;
      17'd58437: data = 8'h19;
      17'd58438: data = 8'h11;
      17'd58439: data = 8'h1f;
      17'd58440: data = 8'hfd;
      17'd58441: data = 8'hfa;
      17'd58442: data = 8'h15;
      17'd58443: data = 8'h06;
      17'd58444: data = 8'h12;
      17'd58445: data = 8'h27;
      17'd58446: data = 8'h24;
      17'd58447: data = 8'h12;
      17'd58448: data = 8'hf6;
      17'd58449: data = 8'he4;
      17'd58450: data = 8'h00;
      17'd58451: data = 8'h04;
      17'd58452: data = 8'h0a;
      17'd58453: data = 8'h29;
      17'd58454: data = 8'h34;
      17'd58455: data = 8'h1c;
      17'd58456: data = 8'h09;
      17'd58457: data = 8'hfa;
      17'd58458: data = 8'hfa;
      17'd58459: data = 8'h06;
      17'd58460: data = 8'hfa;
      17'd58461: data = 8'h02;
      17'd58462: data = 8'hfd;
      17'd58463: data = 8'he3;
      17'd58464: data = 8'h00;
      17'd58465: data = 8'h16;
      17'd58466: data = 8'h1c;
      17'd58467: data = 8'h35;
      17'd58468: data = 8'h29;
      17'd58469: data = 8'h12;
      17'd58470: data = 8'hfd;
      17'd58471: data = 8'hf1;
      17'd58472: data = 8'hf6;
      17'd58473: data = 8'h13;
      17'd58474: data = 8'h1c;
      17'd58475: data = 8'h1b;
      17'd58476: data = 8'h11;
      17'd58477: data = 8'hfa;
      17'd58478: data = 8'hf5;
      17'd58479: data = 8'h05;
      17'd58480: data = 8'h23;
      17'd58481: data = 8'h29;
      17'd58482: data = 8'h1c;
      17'd58483: data = 8'h12;
      17'd58484: data = 8'h00;
      17'd58485: data = 8'hdb;
      17'd58486: data = 8'he3;
      17'd58487: data = 8'h00;
      17'd58488: data = 8'h04;
      17'd58489: data = 8'h09;
      17'd58490: data = 8'h01;
      17'd58491: data = 8'hf4;
      17'd58492: data = 8'hf2;
      17'd58493: data = 8'hed;
      17'd58494: data = 8'hfc;
      17'd58495: data = 8'h09;
      17'd58496: data = 8'hf9;
      17'd58497: data = 8'he5;
      17'd58498: data = 8'hd8;
      17'd58499: data = 8'hcd;
      17'd58500: data = 8'hda;
      17'd58501: data = 8'heb;
      17'd58502: data = 8'hfc;
      17'd58503: data = 8'h04;
      17'd58504: data = 8'hed;
      17'd58505: data = 8'hdc;
      17'd58506: data = 8'hdb;
      17'd58507: data = 8'hda;
      17'd58508: data = 8'hdc;
      17'd58509: data = 8'hf1;
      17'd58510: data = 8'hec;
      17'd58511: data = 8'hde;
      17'd58512: data = 8'hd8;
      17'd58513: data = 8'hd1;
      17'd58514: data = 8'hde;
      17'd58515: data = 8'hf1;
      17'd58516: data = 8'hfe;
      17'd58517: data = 8'h11;
      17'd58518: data = 8'h0a;
      17'd58519: data = 8'hf6;
      17'd58520: data = 8'hf6;
      17'd58521: data = 8'hfd;
      17'd58522: data = 8'hfc;
      17'd58523: data = 8'h02;
      17'd58524: data = 8'h06;
      17'd58525: data = 8'hfd;
      17'd58526: data = 8'hf6;
      17'd58527: data = 8'hf9;
      17'd58528: data = 8'h05;
      17'd58529: data = 8'h1a;
      17'd58530: data = 8'h22;
      17'd58531: data = 8'h23;
      17'd58532: data = 8'h1b;
      17'd58533: data = 8'h0a;
      17'd58534: data = 8'h00;
      17'd58535: data = 8'h02;
      17'd58536: data = 8'h12;
      17'd58537: data = 8'h1b;
      17'd58538: data = 8'h1b;
      17'd58539: data = 8'h19;
      17'd58540: data = 8'h1a;
      17'd58541: data = 8'h12;
      17'd58542: data = 8'h0c;
      17'd58543: data = 8'h19;
      17'd58544: data = 8'h1b;
      17'd58545: data = 8'h12;
      17'd58546: data = 8'h0d;
      17'd58547: data = 8'h06;
      17'd58548: data = 8'h00;
      17'd58549: data = 8'h05;
      17'd58550: data = 8'h0c;
      17'd58551: data = 8'h12;
      17'd58552: data = 8'h13;
      17'd58553: data = 8'h0d;
      17'd58554: data = 8'h0c;
      17'd58555: data = 8'h0a;
      17'd58556: data = 8'h04;
      17'd58557: data = 8'h0a;
      17'd58558: data = 8'h0c;
      17'd58559: data = 8'h05;
      17'd58560: data = 8'hfe;
      17'd58561: data = 8'hf6;
      17'd58562: data = 8'hf6;
      17'd58563: data = 8'hfc;
      17'd58564: data = 8'h04;
      17'd58565: data = 8'h0e;
      17'd58566: data = 8'h16;
      17'd58567: data = 8'h13;
      17'd58568: data = 8'h0e;
      17'd58569: data = 8'h0a;
      17'd58570: data = 8'h05;
      17'd58571: data = 8'h05;
      17'd58572: data = 8'h01;
      17'd58573: data = 8'hf9;
      17'd58574: data = 8'hfa;
      17'd58575: data = 8'hf9;
      17'd58576: data = 8'hf5;
      17'd58577: data = 8'h00;
      17'd58578: data = 8'h04;
      17'd58579: data = 8'h11;
      17'd58580: data = 8'h13;
      17'd58581: data = 8'h0e;
      17'd58582: data = 8'h0c;
      17'd58583: data = 8'h02;
      17'd58584: data = 8'hfc;
      17'd58585: data = 8'hfa;
      17'd58586: data = 8'hfa;
      17'd58587: data = 8'hf9;
      17'd58588: data = 8'hf9;
      17'd58589: data = 8'hf9;
      17'd58590: data = 8'hfe;
      17'd58591: data = 8'h01;
      17'd58592: data = 8'hfd;
      17'd58593: data = 8'hf9;
      17'd58594: data = 8'hf9;
      17'd58595: data = 8'hf5;
      17'd58596: data = 8'hed;
      17'd58597: data = 8'he7;
      17'd58598: data = 8'he3;
      17'd58599: data = 8'he4;
      17'd58600: data = 8'he7;
      17'd58601: data = 8'he7;
      17'd58602: data = 8'he7;
      17'd58603: data = 8'heb;
      17'd58604: data = 8'he7;
      17'd58605: data = 8'he2;
      17'd58606: data = 8'he0;
      17'd58607: data = 8'hdc;
      17'd58608: data = 8'hdb;
      17'd58609: data = 8'hdb;
      17'd58610: data = 8'he0;
      17'd58611: data = 8'he3;
      17'd58612: data = 8'he2;
      17'd58613: data = 8'he2;
      17'd58614: data = 8'he4;
      17'd58615: data = 8'he5;
      17'd58616: data = 8'he7;
      17'd58617: data = 8'hec;
      17'd58618: data = 8'he7;
      17'd58619: data = 8'he3;
      17'd58620: data = 8'hdb;
      17'd58621: data = 8'hd3;
      17'd58622: data = 8'hd8;
      17'd58623: data = 8'hde;
      17'd58624: data = 8'he2;
      17'd58625: data = 8'hed;
      17'd58626: data = 8'hf1;
      17'd58627: data = 8'hef;
      17'd58628: data = 8'hef;
      17'd58629: data = 8'hf4;
      17'd58630: data = 8'hf9;
      17'd58631: data = 8'hf9;
      17'd58632: data = 8'hfa;
      17'd58633: data = 8'hf4;
      17'd58634: data = 8'hf5;
      17'd58635: data = 8'hf1;
      17'd58636: data = 8'hf1;
      17'd58637: data = 8'h00;
      17'd58638: data = 8'h01;
      17'd58639: data = 8'h02;
      17'd58640: data = 8'h0e;
      17'd58641: data = 8'h05;
      17'd58642: data = 8'h02;
      17'd58643: data = 8'h0e;
      17'd58644: data = 8'h0c;
      17'd58645: data = 8'h15;
      17'd58646: data = 8'h1a;
      17'd58647: data = 8'h0c;
      17'd58648: data = 8'h09;
      17'd58649: data = 8'h0c;
      17'd58650: data = 8'h05;
      17'd58651: data = 8'h15;
      17'd58652: data = 8'h12;
      17'd58653: data = 8'h16;
      17'd58654: data = 8'h1b;
      17'd58655: data = 8'h13;
      17'd58656: data = 8'h0a;
      17'd58657: data = 8'h12;
      17'd58658: data = 8'h04;
      17'd58659: data = 8'h06;
      17'd58660: data = 8'h1c;
      17'd58661: data = 8'h02;
      17'd58662: data = 8'h12;
      17'd58663: data = 8'h1a;
      17'd58664: data = 8'h01;
      17'd58665: data = 8'h16;
      17'd58666: data = 8'h1f;
      17'd58667: data = 8'h06;
      17'd58668: data = 8'h00;
      17'd58669: data = 8'h11;
      17'd58670: data = 8'h00;
      17'd58671: data = 8'hfa;
      17'd58672: data = 8'h05;
      17'd58673: data = 8'h0d;
      17'd58674: data = 8'h05;
      17'd58675: data = 8'h04;
      17'd58676: data = 8'h16;
      17'd58677: data = 8'h1e;
      17'd58678: data = 8'h22;
      17'd58679: data = 8'h23;
      17'd58680: data = 8'h1b;
      17'd58681: data = 8'h02;
      17'd58682: data = 8'h00;
      17'd58683: data = 8'he4;
      17'd58684: data = 8'hce;
      17'd58685: data = 8'hfd;
      17'd58686: data = 8'h09;
      17'd58687: data = 8'h02;
      17'd58688: data = 8'h27;
      17'd58689: data = 8'h36;
      17'd58690: data = 8'h15;
      17'd58691: data = 8'h0a;
      17'd58692: data = 8'h00;
      17'd58693: data = 8'h04;
      17'd58694: data = 8'h13;
      17'd58695: data = 8'hfe;
      17'd58696: data = 8'hed;
      17'd58697: data = 8'h13;
      17'd58698: data = 8'h1b;
      17'd58699: data = 8'h13;
      17'd58700: data = 8'h23;
      17'd58701: data = 8'h2b;
      17'd58702: data = 8'h2b;
      17'd58703: data = 8'h13;
      17'd58704: data = 8'h00;
      17'd58705: data = 8'hfa;
      17'd58706: data = 8'h00;
      17'd58707: data = 8'h01;
      17'd58708: data = 8'h0d;
      17'd58709: data = 8'h05;
      17'd58710: data = 8'h04;
      17'd58711: data = 8'h01;
      17'd58712: data = 8'hf2;
      17'd58713: data = 8'h09;
      17'd58714: data = 8'h0d;
      17'd58715: data = 8'hfc;
      17'd58716: data = 8'h01;
      17'd58717: data = 8'h02;
      17'd58718: data = 8'he0;
      17'd58719: data = 8'he2;
      17'd58720: data = 8'he5;
      17'd58721: data = 8'he9;
      17'd58722: data = 8'h01;
      17'd58723: data = 8'hfd;
      17'd58724: data = 8'hf4;
      17'd58725: data = 8'hfd;
      17'd58726: data = 8'hf5;
      17'd58727: data = 8'he9;
      17'd58728: data = 8'hed;
      17'd58729: data = 8'he0;
      17'd58730: data = 8'he0;
      17'd58731: data = 8'hd8;
      17'd58732: data = 8'hcd;
      17'd58733: data = 8'hde;
      17'd58734: data = 8'he5;
      17'd58735: data = 8'heb;
      17'd58736: data = 8'hfe;
      17'd58737: data = 8'hfc;
      17'd58738: data = 8'hef;
      17'd58739: data = 8'hf2;
      17'd58740: data = 8'he9;
      17'd58741: data = 8'he9;
      17'd58742: data = 8'hf5;
      17'd58743: data = 8'hf1;
      17'd58744: data = 8'hf4;
      17'd58745: data = 8'h02;
      17'd58746: data = 8'hfe;
      17'd58747: data = 8'h04;
      17'd58748: data = 8'h0a;
      17'd58749: data = 8'h0a;
      17'd58750: data = 8'h11;
      17'd58751: data = 8'h0c;
      17'd58752: data = 8'h00;
      17'd58753: data = 8'hfd;
      17'd58754: data = 8'h01;
      17'd58755: data = 8'h01;
      17'd58756: data = 8'h0a;
      17'd58757: data = 8'h0e;
      17'd58758: data = 8'h11;
      17'd58759: data = 8'h19;
      17'd58760: data = 8'h13;
      17'd58761: data = 8'h11;
      17'd58762: data = 8'h16;
      17'd58763: data = 8'h13;
      17'd58764: data = 8'h0d;
      17'd58765: data = 8'h0a;
      17'd58766: data = 8'h05;
      17'd58767: data = 8'h04;
      17'd58768: data = 8'h09;
      17'd58769: data = 8'h0d;
      17'd58770: data = 8'h16;
      17'd58771: data = 8'h1c;
      17'd58772: data = 8'h19;
      17'd58773: data = 8'h16;
      17'd58774: data = 8'h12;
      17'd58775: data = 8'h04;
      17'd58776: data = 8'h05;
      17'd58777: data = 8'h02;
      17'd58778: data = 8'hfe;
      17'd58779: data = 8'h02;
      17'd58780: data = 8'h01;
      17'd58781: data = 8'h04;
      17'd58782: data = 8'h0d;
      17'd58783: data = 8'h0e;
      17'd58784: data = 8'h0a;
      17'd58785: data = 8'h0a;
      17'd58786: data = 8'h05;
      17'd58787: data = 8'h00;
      17'd58788: data = 8'h02;
      17'd58789: data = 8'h02;
      17'd58790: data = 8'h06;
      17'd58791: data = 8'h0d;
      17'd58792: data = 8'h09;
      17'd58793: data = 8'h0c;
      17'd58794: data = 8'h0d;
      17'd58795: data = 8'h06;
      17'd58796: data = 8'h06;
      17'd58797: data = 8'h04;
      17'd58798: data = 8'h01;
      17'd58799: data = 8'h00;
      17'd58800: data = 8'hfd;
      17'd58801: data = 8'hfe;
      17'd58802: data = 8'h04;
      17'd58803: data = 8'h02;
      17'd58804: data = 8'h02;
      17'd58805: data = 8'h05;
      17'd58806: data = 8'h02;
      17'd58807: data = 8'h01;
      17'd58808: data = 8'h01;
      17'd58809: data = 8'hfd;
      17'd58810: data = 8'h01;
      17'd58811: data = 8'h00;
      17'd58812: data = 8'hf9;
      17'd58813: data = 8'hfa;
      17'd58814: data = 8'hf6;
      17'd58815: data = 8'hf5;
      17'd58816: data = 8'hfd;
      17'd58817: data = 8'hfa;
      17'd58818: data = 8'hf9;
      17'd58819: data = 8'hf9;
      17'd58820: data = 8'hf4;
      17'd58821: data = 8'hf1;
      17'd58822: data = 8'heb;
      17'd58823: data = 8'he7;
      17'd58824: data = 8'he7;
      17'd58825: data = 8'he5;
      17'd58826: data = 8'he4;
      17'd58827: data = 8'he5;
      17'd58828: data = 8'he7;
      17'd58829: data = 8'he5;
      17'd58830: data = 8'he9;
      17'd58831: data = 8'he4;
      17'd58832: data = 8'hde;
      17'd58833: data = 8'he2;
      17'd58834: data = 8'he2;
      17'd58835: data = 8'he2;
      17'd58836: data = 8'he3;
      17'd58837: data = 8'he4;
      17'd58838: data = 8'he5;
      17'd58839: data = 8'he5;
      17'd58840: data = 8'he2;
      17'd58841: data = 8'he2;
      17'd58842: data = 8'he4;
      17'd58843: data = 8'he0;
      17'd58844: data = 8'he3;
      17'd58845: data = 8'he2;
      17'd58846: data = 8'hdc;
      17'd58847: data = 8'he3;
      17'd58848: data = 8'he2;
      17'd58849: data = 8'he5;
      17'd58850: data = 8'hed;
      17'd58851: data = 8'hed;
      17'd58852: data = 8'hf1;
      17'd58853: data = 8'hf5;
      17'd58854: data = 8'hf4;
      17'd58855: data = 8'hf1;
      17'd58856: data = 8'hf5;
      17'd58857: data = 8'hf4;
      17'd58858: data = 8'hf4;
      17'd58859: data = 8'hf6;
      17'd58860: data = 8'hfa;
      17'd58861: data = 8'hfc;
      17'd58862: data = 8'hfd;
      17'd58863: data = 8'h04;
      17'd58864: data = 8'h06;
      17'd58865: data = 8'h09;
      17'd58866: data = 8'h0a;
      17'd58867: data = 8'h0a;
      17'd58868: data = 8'h04;
      17'd58869: data = 8'h09;
      17'd58870: data = 8'h0e;
      17'd58871: data = 8'h06;
      17'd58872: data = 8'h0c;
      17'd58873: data = 8'h0c;
      17'd58874: data = 8'h0e;
      17'd58875: data = 8'h0c;
      17'd58876: data = 8'h0a;
      17'd58877: data = 8'h12;
      17'd58878: data = 8'h0c;
      17'd58879: data = 8'h13;
      17'd58880: data = 8'h12;
      17'd58881: data = 8'h12;
      17'd58882: data = 8'h0c;
      17'd58883: data = 8'h06;
      17'd58884: data = 8'h16;
      17'd58885: data = 8'h15;
      17'd58886: data = 8'h15;
      17'd58887: data = 8'h0a;
      17'd58888: data = 8'h19;
      17'd58889: data = 8'h11;
      17'd58890: data = 8'h01;
      17'd58891: data = 8'h12;
      17'd58892: data = 8'h00;
      17'd58893: data = 8'h09;
      17'd58894: data = 8'h19;
      17'd58895: data = 8'h04;
      17'd58896: data = 8'h12;
      17'd58897: data = 8'h15;
      17'd58898: data = 8'hfc;
      17'd58899: data = 8'h1a;
      17'd58900: data = 8'h16;
      17'd58901: data = 8'h13;
      17'd58902: data = 8'h09;
      17'd58903: data = 8'h05;
      17'd58904: data = 8'h06;
      17'd58905: data = 8'hf9;
      17'd58906: data = 8'h06;
      17'd58907: data = 8'h19;
      17'd58908: data = 8'h35;
      17'd58909: data = 8'h29;
      17'd58910: data = 8'h13;
      17'd58911: data = 8'h0e;
      17'd58912: data = 8'he0;
      17'd58913: data = 8'hd8;
      17'd58914: data = 8'hfd;
      17'd58915: data = 8'hf9;
      17'd58916: data = 8'h11;
      17'd58917: data = 8'h27;
      17'd58918: data = 8'h0e;
      17'd58919: data = 8'h0d;
      17'd58920: data = 8'h05;
      17'd58921: data = 8'h06;
      17'd58922: data = 8'h0c;
      17'd58923: data = 8'h02;
      17'd58924: data = 8'hf4;
      17'd58925: data = 8'he7;
      17'd58926: data = 8'hf9;
      17'd58927: data = 8'hf6;
      17'd58928: data = 8'h24;
      17'd58929: data = 8'h2d;
      17'd58930: data = 8'h1f;
      17'd58931: data = 8'h27;
      17'd58932: data = 8'h01;
      17'd58933: data = 8'hec;
      17'd58934: data = 8'hec;
      17'd58935: data = 8'hfc;
      17'd58936: data = 8'h0a;
      17'd58937: data = 8'h0d;
      17'd58938: data = 8'h0a;
      17'd58939: data = 8'h02;
      17'd58940: data = 8'h01;
      17'd58941: data = 8'hf5;
      17'd58942: data = 8'hfc;
      17'd58943: data = 8'h09;
      17'd58944: data = 8'hef;
      17'd58945: data = 8'hf9;
      17'd58946: data = 8'hf6;
      17'd58947: data = 8'he2;
      17'd58948: data = 8'hf5;
      17'd58949: data = 8'hfe;
      17'd58950: data = 8'hfe;
      17'd58951: data = 8'h04;
      17'd58952: data = 8'hfe;
      17'd58953: data = 8'hf1;
      17'd58954: data = 8'he9;
      17'd58955: data = 8'heb;
      17'd58956: data = 8'he7;
      17'd58957: data = 8'hf6;
      17'd58958: data = 8'hef;
      17'd58959: data = 8'heb;
      17'd58960: data = 8'hf1;
      17'd58961: data = 8'hde;
      17'd58962: data = 8'he5;
      17'd58963: data = 8'hf1;
      17'd58964: data = 8'hf1;
      17'd58965: data = 8'hf5;
      17'd58966: data = 8'hed;
      17'd58967: data = 8'he9;
      17'd58968: data = 8'he4;
      17'd58969: data = 8'he0;
      17'd58970: data = 8'he9;
      17'd58971: data = 8'hf5;
      17'd58972: data = 8'hfa;
      17'd58973: data = 8'hfd;
      17'd58974: data = 8'h05;
      17'd58975: data = 8'h00;
      17'd58976: data = 8'h00;
      17'd58977: data = 8'h0a;
      17'd58978: data = 8'h0a;
      17'd58979: data = 8'h0a;
      17'd58980: data = 8'h05;
      17'd58981: data = 8'hfe;
      17'd58982: data = 8'hfe;
      17'd58983: data = 8'h00;
      17'd58984: data = 8'h09;
      17'd58985: data = 8'h15;
      17'd58986: data = 8'h19;
      17'd58987: data = 8'h16;
      17'd58988: data = 8'h11;
      17'd58989: data = 8'h05;
      17'd58990: data = 8'h02;
      17'd58991: data = 8'h0a;
      17'd58992: data = 8'h0e;
      17'd58993: data = 8'h11;
      17'd58994: data = 8'h1a;
      17'd58995: data = 8'h19;
      17'd58996: data = 8'h19;
      17'd58997: data = 8'h1a;
      17'd58998: data = 8'h19;
      17'd58999: data = 8'h1a;
      17'd59000: data = 8'h19;
      17'd59001: data = 8'h13;
      17'd59002: data = 8'h0d;
      17'd59003: data = 8'h09;
      17'd59004: data = 8'h06;
      17'd59005: data = 8'h0c;
      17'd59006: data = 8'h12;
      17'd59007: data = 8'h0e;
      17'd59008: data = 8'h11;
      17'd59009: data = 8'h0e;
      17'd59010: data = 8'h06;
      17'd59011: data = 8'h05;
      17'd59012: data = 8'h05;
      17'd59013: data = 8'h04;
      17'd59014: data = 8'h05;
      17'd59015: data = 8'h04;
      17'd59016: data = 8'h01;
      17'd59017: data = 8'h00;
      17'd59018: data = 8'hfe;
      17'd59019: data = 8'h01;
      17'd59020: data = 8'h02;
      17'd59021: data = 8'h01;
      17'd59022: data = 8'h02;
      17'd59023: data = 8'h02;
      17'd59024: data = 8'h01;
      17'd59025: data = 8'h02;
      17'd59026: data = 8'h04;
      17'd59027: data = 8'h00;
      17'd59028: data = 8'h01;
      17'd59029: data = 8'h01;
      17'd59030: data = 8'hfe;
      17'd59031: data = 8'h00;
      17'd59032: data = 8'h02;
      17'd59033: data = 8'h00;
      17'd59034: data = 8'hfd;
      17'd59035: data = 8'hfd;
      17'd59036: data = 8'hfc;
      17'd59037: data = 8'hfa;
      17'd59038: data = 8'hfd;
      17'd59039: data = 8'h00;
      17'd59040: data = 8'hfd;
      17'd59041: data = 8'h00;
      17'd59042: data = 8'h01;
      17'd59043: data = 8'h00;
      17'd59044: data = 8'h00;
      17'd59045: data = 8'hfe;
      17'd59046: data = 8'hf9;
      17'd59047: data = 8'hf5;
      17'd59048: data = 8'hf2;
      17'd59049: data = 8'hef;
      17'd59050: data = 8'hf1;
      17'd59051: data = 8'hf1;
      17'd59052: data = 8'hf1;
      17'd59053: data = 8'hf2;
      17'd59054: data = 8'hef;
      17'd59055: data = 8'hed;
      17'd59056: data = 8'he9;
      17'd59057: data = 8'he4;
      17'd59058: data = 8'he5;
      17'd59059: data = 8'he4;
      17'd59060: data = 8'he2;
      17'd59061: data = 8'he4;
      17'd59062: data = 8'he2;
      17'd59063: data = 8'hde;
      17'd59064: data = 8'he5;
      17'd59065: data = 8'he4;
      17'd59066: data = 8'he2;
      17'd59067: data = 8'he4;
      17'd59068: data = 8'he0;
      17'd59069: data = 8'hde;
      17'd59070: data = 8'hde;
      17'd59071: data = 8'he2;
      17'd59072: data = 8'he7;
      17'd59073: data = 8'hed;
      17'd59074: data = 8'hec;
      17'd59075: data = 8'hec;
      17'd59076: data = 8'he9;
      17'd59077: data = 8'he5;
      17'd59078: data = 8'he5;
      17'd59079: data = 8'he9;
      17'd59080: data = 8'hec;
      17'd59081: data = 8'hef;
      17'd59082: data = 8'hed;
      17'd59083: data = 8'hef;
      17'd59084: data = 8'hf4;
      17'd59085: data = 8'hf9;
      17'd59086: data = 8'hfd;
      17'd59087: data = 8'h01;
      17'd59088: data = 8'h01;
      17'd59089: data = 8'h01;
      17'd59090: data = 8'hfe;
      17'd59091: data = 8'hfe;
      17'd59092: data = 8'h04;
      17'd59093: data = 8'h0a;
      17'd59094: data = 8'h0a;
      17'd59095: data = 8'h06;
      17'd59096: data = 8'h09;
      17'd59097: data = 8'h06;
      17'd59098: data = 8'h04;
      17'd59099: data = 8'h0c;
      17'd59100: data = 8'h0d;
      17'd59101: data = 8'h0c;
      17'd59102: data = 8'h11;
      17'd59103: data = 8'h11;
      17'd59104: data = 8'h0a;
      17'd59105: data = 8'h0a;
      17'd59106: data = 8'h0a;
      17'd59107: data = 8'h0c;
      17'd59108: data = 8'h13;
      17'd59109: data = 8'h09;
      17'd59110: data = 8'h05;
      17'd59111: data = 8'h09;
      17'd59112: data = 8'h06;
      17'd59113: data = 8'h0a;
      17'd59114: data = 8'h0c;
      17'd59115: data = 8'h05;
      17'd59116: data = 8'h09;
      17'd59117: data = 8'h0a;
      17'd59118: data = 8'h05;
      17'd59119: data = 8'h05;
      17'd59120: data = 8'h0e;
      17'd59121: data = 8'h09;
      17'd59122: data = 8'h0d;
      17'd59123: data = 8'h0d;
      17'd59124: data = 8'h05;
      17'd59125: data = 8'h06;
      17'd59126: data = 8'h02;
      17'd59127: data = 8'h0d;
      17'd59128: data = 8'h02;
      17'd59129: data = 8'h06;
      17'd59130: data = 8'h0c;
      17'd59131: data = 8'h02;
      17'd59132: data = 8'h06;
      17'd59133: data = 8'h0d;
      17'd59134: data = 8'h06;
      17'd59135: data = 8'h06;
      17'd59136: data = 8'h0d;
      17'd59137: data = 8'h09;
      17'd59138: data = 8'h05;
      17'd59139: data = 8'h0d;
      17'd59140: data = 8'h0a;
      17'd59141: data = 8'h0d;
      17'd59142: data = 8'h12;
      17'd59143: data = 8'h0e;
      17'd59144: data = 8'h02;
      17'd59145: data = 8'hfe;
      17'd59146: data = 8'hf9;
      17'd59147: data = 8'h00;
      17'd59148: data = 8'h00;
      17'd59149: data = 8'hfe;
      17'd59150: data = 8'h0a;
      17'd59151: data = 8'h0d;
      17'd59152: data = 8'h0c;
      17'd59153: data = 8'h01;
      17'd59154: data = 8'hfc;
      17'd59155: data = 8'hf5;
      17'd59156: data = 8'hf9;
      17'd59157: data = 8'hf6;
      17'd59158: data = 8'hf2;
      17'd59159: data = 8'hf5;
      17'd59160: data = 8'h02;
      17'd59161: data = 8'h0a;
      17'd59162: data = 8'h0c;
      17'd59163: data = 8'h04;
      17'd59164: data = 8'h04;
      17'd59165: data = 8'h05;
      17'd59166: data = 8'hfc;
      17'd59167: data = 8'hf9;
      17'd59168: data = 8'hfa;
      17'd59169: data = 8'h00;
      17'd59170: data = 8'h06;
      17'd59171: data = 8'h0c;
      17'd59172: data = 8'h06;
      17'd59173: data = 8'h01;
      17'd59174: data = 8'h01;
      17'd59175: data = 8'hfd;
      17'd59176: data = 8'hfc;
      17'd59177: data = 8'hf6;
      17'd59178: data = 8'hfa;
      17'd59179: data = 8'h00;
      17'd59180: data = 8'hfe;
      17'd59181: data = 8'h01;
      17'd59182: data = 8'h01;
      17'd59183: data = 8'h05;
      17'd59184: data = 8'h0c;
      17'd59185: data = 8'h0a;
      17'd59186: data = 8'h01;
      17'd59187: data = 8'h01;
      17'd59188: data = 8'hfe;
      17'd59189: data = 8'hf9;
      17'd59190: data = 8'hf9;
      17'd59191: data = 8'hf9;
      17'd59192: data = 8'hfc;
      17'd59193: data = 8'hfe;
      17'd59194: data = 8'h00;
      17'd59195: data = 8'hfe;
      17'd59196: data = 8'hfa;
      17'd59197: data = 8'hf6;
      17'd59198: data = 8'hf6;
      17'd59199: data = 8'hf4;
      17'd59200: data = 8'hf1;
      17'd59201: data = 8'hf1;
      17'd59202: data = 8'hf4;
      17'd59203: data = 8'hf9;
      17'd59204: data = 8'hfc;
      17'd59205: data = 8'hfc;
      17'd59206: data = 8'hfc;
      17'd59207: data = 8'hfd;
      17'd59208: data = 8'hf9;
      17'd59209: data = 8'hf9;
      17'd59210: data = 8'hf6;
      17'd59211: data = 8'hf6;
      17'd59212: data = 8'hfc;
      17'd59213: data = 8'h00;
      17'd59214: data = 8'h04;
      17'd59215: data = 8'h05;
      17'd59216: data = 8'h0a;
      17'd59217: data = 8'h06;
      17'd59218: data = 8'h05;
      17'd59219: data = 8'h05;
      17'd59220: data = 8'h04;
      17'd59221: data = 8'h04;
      17'd59222: data = 8'h02;
      17'd59223: data = 8'h04;
      17'd59224: data = 8'h01;
      17'd59225: data = 8'h04;
      17'd59226: data = 8'h05;
      17'd59227: data = 8'h05;
      17'd59228: data = 8'h0a;
      17'd59229: data = 8'h0c;
      17'd59230: data = 8'h0c;
      17'd59231: data = 8'h0a;
      17'd59232: data = 8'h09;
      17'd59233: data = 8'h0a;
      17'd59234: data = 8'h0c;
      17'd59235: data = 8'h0c;
      17'd59236: data = 8'h0a;
      17'd59237: data = 8'h09;
      17'd59238: data = 8'h06;
      17'd59239: data = 8'h05;
      17'd59240: data = 8'h04;
      17'd59241: data = 8'h02;
      17'd59242: data = 8'h01;
      17'd59243: data = 8'h02;
      17'd59244: data = 8'h01;
      17'd59245: data = 8'h01;
      17'd59246: data = 8'hfe;
      17'd59247: data = 8'hfe;
      17'd59248: data = 8'hfe;
      17'd59249: data = 8'hfe;
      17'd59250: data = 8'hfd;
      17'd59251: data = 8'hfc;
      17'd59252: data = 8'hfa;
      17'd59253: data = 8'hfd;
      17'd59254: data = 8'hfd;
      17'd59255: data = 8'hfe;
      17'd59256: data = 8'h00;
      17'd59257: data = 8'hfc;
      17'd59258: data = 8'hfd;
      17'd59259: data = 8'hfe;
      17'd59260: data = 8'hfd;
      17'd59261: data = 8'hfd;
      17'd59262: data = 8'hfd;
      17'd59263: data = 8'hfd;
      17'd59264: data = 8'hfe;
      17'd59265: data = 8'hfd;
      17'd59266: data = 8'hfc;
      17'd59267: data = 8'hfe;
      17'd59268: data = 8'hfd;
      17'd59269: data = 8'hfd;
      17'd59270: data = 8'hfd;
      17'd59271: data = 8'hfa;
      17'd59272: data = 8'hfa;
      17'd59273: data = 8'hfa;
      17'd59274: data = 8'hf9;
      17'd59275: data = 8'hfc;
      17'd59276: data = 8'hfd;
      17'd59277: data = 8'hfe;
      17'd59278: data = 8'h02;
      17'd59279: data = 8'hfe;
      17'd59280: data = 8'hfc;
      17'd59281: data = 8'hfd;
      17'd59282: data = 8'hfc;
      17'd59283: data = 8'hf9;
      17'd59284: data = 8'hf6;
      17'd59285: data = 8'hf9;
      17'd59286: data = 8'hf6;
      17'd59287: data = 8'hf6;
      17'd59288: data = 8'hf5;
      17'd59289: data = 8'hf5;
      17'd59290: data = 8'hf5;
      17'd59291: data = 8'hf2;
      17'd59292: data = 8'hf2;
      17'd59293: data = 8'hef;
      17'd59294: data = 8'hed;
      17'd59295: data = 8'hec;
      17'd59296: data = 8'heb;
      17'd59297: data = 8'hed;
      17'd59298: data = 8'hed;
      17'd59299: data = 8'hed;
      17'd59300: data = 8'hed;
      17'd59301: data = 8'hec;
      17'd59302: data = 8'heb;
      17'd59303: data = 8'he9;
      17'd59304: data = 8'he9;
      17'd59305: data = 8'hec;
      17'd59306: data = 8'hed;
      17'd59307: data = 8'hed;
      17'd59308: data = 8'hf1;
      17'd59309: data = 8'hef;
      17'd59310: data = 8'hec;
      17'd59311: data = 8'hec;
      17'd59312: data = 8'hed;
      17'd59313: data = 8'hed;
      17'd59314: data = 8'hef;
      17'd59315: data = 8'hef;
      17'd59316: data = 8'hef;
      17'd59317: data = 8'hf1;
      17'd59318: data = 8'hf4;
      17'd59319: data = 8'hf6;
      17'd59320: data = 8'hf9;
      17'd59321: data = 8'hf9;
      17'd59322: data = 8'hf9;
      17'd59323: data = 8'hf5;
      17'd59324: data = 8'hf6;
      17'd59325: data = 8'hfe;
      17'd59326: data = 8'hfd;
      17'd59327: data = 8'h00;
      17'd59328: data = 8'h02;
      17'd59329: data = 8'h01;
      17'd59330: data = 8'hfe;
      17'd59331: data = 8'hfe;
      17'd59332: data = 8'h00;
      17'd59333: data = 8'h02;
      17'd59334: data = 8'h04;
      17'd59335: data = 8'h04;
      17'd59336: data = 8'h04;
      17'd59337: data = 8'h05;
      17'd59338: data = 8'h05;
      17'd59339: data = 8'h04;
      17'd59340: data = 8'h04;
      17'd59341: data = 8'h06;
      17'd59342: data = 8'h09;
      17'd59343: data = 8'h09;
      17'd59344: data = 8'h06;
      17'd59345: data = 8'h06;
      17'd59346: data = 8'h0c;
      17'd59347: data = 8'h0d;
      17'd59348: data = 8'h0a;
      17'd59349: data = 8'h06;
      17'd59350: data = 8'h06;
      17'd59351: data = 8'h06;
      17'd59352: data = 8'h06;
      17'd59353: data = 8'h09;
      17'd59354: data = 8'h06;
      17'd59355: data = 8'h09;
      17'd59356: data = 8'h0c;
      17'd59357: data = 8'h0c;
      17'd59358: data = 8'h06;
      17'd59359: data = 8'h05;
      17'd59360: data = 8'h0a;
      17'd59361: data = 8'h0a;
      17'd59362: data = 8'h0c;
      17'd59363: data = 8'h09;
      17'd59364: data = 8'h04;
      17'd59365: data = 8'h05;
      17'd59366: data = 8'h09;
      17'd59367: data = 8'h06;
      17'd59368: data = 8'h05;
      17'd59369: data = 8'h0a;
      17'd59370: data = 8'h0c;
      17'd59371: data = 8'h0a;
      17'd59372: data = 8'h0a;
      17'd59373: data = 8'h0c;
      17'd59374: data = 8'h0d;
      17'd59375: data = 8'h0d;
      17'd59376: data = 8'h0c;
      17'd59377: data = 8'h0a;
      17'd59378: data = 8'h0e;
      17'd59379: data = 8'h0e;
      17'd59380: data = 8'h05;
      17'd59381: data = 8'h02;
      17'd59382: data = 8'h02;
      17'd59383: data = 8'hfd;
      17'd59384: data = 8'hf9;
      17'd59385: data = 8'hfe;
      17'd59386: data = 8'h05;
      17'd59387: data = 8'h06;
      17'd59388: data = 8'h04;
      17'd59389: data = 8'h06;
      17'd59390: data = 8'h0a;
      17'd59391: data = 8'h05;
      17'd59392: data = 8'hfd;
      17'd59393: data = 8'hf9;
      17'd59394: data = 8'h00;
      17'd59395: data = 8'h01;
      17'd59396: data = 8'hfd;
      17'd59397: data = 8'h00;
      17'd59398: data = 8'h05;
      17'd59399: data = 8'h0d;
      17'd59400: data = 8'h0d;
      17'd59401: data = 8'h06;
      17'd59402: data = 8'h06;
      17'd59403: data = 8'h06;
      17'd59404: data = 8'h05;
      17'd59405: data = 8'h04;
      17'd59406: data = 8'h02;
      17'd59407: data = 8'h01;
      17'd59408: data = 8'h02;
      17'd59409: data = 8'h09;
      17'd59410: data = 8'h06;
      17'd59411: data = 8'h02;
      17'd59412: data = 8'h01;
      17'd59413: data = 8'h02;
      17'd59414: data = 8'h05;
      17'd59415: data = 8'hfe;
      17'd59416: data = 8'hfd;
      17'd59417: data = 8'h02;
      17'd59418: data = 8'h0a;
      17'd59419: data = 8'h0c;
      17'd59420: data = 8'h09;
      17'd59421: data = 8'h11;
      17'd59422: data = 8'h0e;
      17'd59423: data = 8'h09;
      17'd59424: data = 8'h05;
      17'd59425: data = 8'h01;
      17'd59426: data = 8'hfe;
      17'd59427: data = 8'hfd;
      17'd59428: data = 8'hfc;
      17'd59429: data = 8'hfa;
      17'd59430: data = 8'hfd;
      17'd59431: data = 8'hfc;
      17'd59432: data = 8'hf9;
      17'd59433: data = 8'hfa;
      17'd59434: data = 8'hfc;
      17'd59435: data = 8'hf5;
      17'd59436: data = 8'hf4;
      17'd59437: data = 8'hfa;
      17'd59438: data = 8'hf9;
      17'd59439: data = 8'hf6;
      17'd59440: data = 8'hfc;
      17'd59441: data = 8'hfe;
      17'd59442: data = 8'hfd;
      17'd59443: data = 8'hf9;
      17'd59444: data = 8'hf9;
      17'd59445: data = 8'hf5;
      17'd59446: data = 8'hf5;
      17'd59447: data = 8'hf5;
      17'd59448: data = 8'hf9;
      17'd59449: data = 8'hfd;
      17'd59450: data = 8'h02;
      17'd59451: data = 8'h05;
      17'd59452: data = 8'h01;
      17'd59453: data = 8'h04;
      17'd59454: data = 8'h01;
      17'd59455: data = 8'hfe;
      17'd59456: data = 8'hf9;
      17'd59457: data = 8'hfa;
      17'd59458: data = 8'hfd;
      17'd59459: data = 8'hfc;
      17'd59460: data = 8'hfe;
      17'd59461: data = 8'hfe;
      17'd59462: data = 8'h04;
      17'd59463: data = 8'h06;
      17'd59464: data = 8'h04;
      17'd59465: data = 8'h04;
      17'd59466: data = 8'h04;
      17'd59467: data = 8'h05;
      17'd59468: data = 8'h05;
      17'd59469: data = 8'h05;
      17'd59470: data = 8'h0a;
      17'd59471: data = 8'h0c;
      17'd59472: data = 8'h0e;
      17'd59473: data = 8'h0d;
      17'd59474: data = 8'h0a;
      17'd59475: data = 8'h02;
      17'd59476: data = 8'h00;
      17'd59477: data = 8'h00;
      17'd59478: data = 8'h00;
      17'd59479: data = 8'h01;
      17'd59480: data = 8'h02;
      17'd59481: data = 8'h05;
      17'd59482: data = 8'h06;
      17'd59483: data = 8'h09;
      17'd59484: data = 8'h05;
      17'd59485: data = 8'h05;
      17'd59486: data = 8'h02;
      17'd59487: data = 8'h00;
      17'd59488: data = 8'hfc;
      17'd59489: data = 8'hfe;
      17'd59490: data = 8'hfe;
      17'd59491: data = 8'h00;
      17'd59492: data = 8'h02;
      17'd59493: data = 8'h01;
      17'd59494: data = 8'h01;
      17'd59495: data = 8'h00;
      17'd59496: data = 8'hfd;
      17'd59497: data = 8'hfc;
      17'd59498: data = 8'hfd;
      17'd59499: data = 8'h00;
      17'd59500: data = 8'h00;
      17'd59501: data = 8'hfe;
      17'd59502: data = 8'h00;
      17'd59503: data = 8'hfe;
      17'd59504: data = 8'hfe;
      17'd59505: data = 8'hfc;
      17'd59506: data = 8'hfa;
      17'd59507: data = 8'hfa;
      17'd59508: data = 8'hfa;
      17'd59509: data = 8'hf9;
      17'd59510: data = 8'hf6;
      17'd59511: data = 8'hfc;
      17'd59512: data = 8'hfc;
      17'd59513: data = 8'hfd;
      17'd59514: data = 8'hfe;
      17'd59515: data = 8'hfe;
      17'd59516: data = 8'hfd;
      17'd59517: data = 8'hfa;
      17'd59518: data = 8'hfa;
      17'd59519: data = 8'hf9;
      17'd59520: data = 8'hf6;
      17'd59521: data = 8'hf5;
      17'd59522: data = 8'hf5;
      17'd59523: data = 8'hf5;
      17'd59524: data = 8'hf1;
      17'd59525: data = 8'hf1;
      17'd59526: data = 8'hef;
      17'd59527: data = 8'hef;
      17'd59528: data = 8'hf1;
      17'd59529: data = 8'hf1;
      17'd59530: data = 8'hef;
      17'd59531: data = 8'hed;
      17'd59532: data = 8'hec;
      17'd59533: data = 8'hef;
      17'd59534: data = 8'hef;
      17'd59535: data = 8'hf1;
      17'd59536: data = 8'hec;
      17'd59537: data = 8'hed;
      17'd59538: data = 8'hec;
      17'd59539: data = 8'he9;
      17'd59540: data = 8'heb;
      17'd59541: data = 8'heb;
      17'd59542: data = 8'hec;
      17'd59543: data = 8'hec;
      17'd59544: data = 8'hec;
      17'd59545: data = 8'hec;
      17'd59546: data = 8'hed;
      17'd59547: data = 8'hef;
      17'd59548: data = 8'hed;
      17'd59549: data = 8'hed;
      17'd59550: data = 8'hed;
      17'd59551: data = 8'hed;
      17'd59552: data = 8'heb;
      17'd59553: data = 8'hec;
      17'd59554: data = 8'hec;
      17'd59555: data = 8'hef;
      17'd59556: data = 8'hf2;
      17'd59557: data = 8'hf2;
      17'd59558: data = 8'hf2;
      17'd59559: data = 8'hf4;
      17'd59560: data = 8'hf9;
      17'd59561: data = 8'hfa;
      17'd59562: data = 8'hfc;
      17'd59563: data = 8'h01;
      17'd59564: data = 8'h00;
      17'd59565: data = 8'h00;
      17'd59566: data = 8'h01;
      17'd59567: data = 8'h01;
      17'd59568: data = 8'h00;
      17'd59569: data = 8'h01;
      17'd59570: data = 8'h02;
      17'd59571: data = 8'h02;
      17'd59572: data = 8'h01;
      17'd59573: data = 8'h01;
      17'd59574: data = 8'h02;
      17'd59575: data = 8'h05;
      17'd59576: data = 8'h09;
      17'd59577: data = 8'h06;
      17'd59578: data = 8'h09;
      17'd59579: data = 8'h0c;
      17'd59580: data = 8'h0a;
      17'd59581: data = 8'h0a;
      17'd59582: data = 8'h0a;
      17'd59583: data = 8'h09;
      17'd59584: data = 8'h0a;
      17'd59585: data = 8'h0c;
      17'd59586: data = 8'h0a;
      17'd59587: data = 8'h09;
      17'd59588: data = 8'h0a;
      17'd59589: data = 8'h0a;
      17'd59590: data = 8'h0d;
      17'd59591: data = 8'h0d;
      17'd59592: data = 8'h0c;
      17'd59593: data = 8'h0c;
      17'd59594: data = 8'h0d;
      17'd59595: data = 8'h0d;
      17'd59596: data = 8'h0e;
      17'd59597: data = 8'h11;
      17'd59598: data = 8'h0c;
      17'd59599: data = 8'h0a;
      17'd59600: data = 8'h06;
      17'd59601: data = 8'h04;
      17'd59602: data = 8'h02;
      17'd59603: data = 8'h05;
      17'd59604: data = 8'h09;
      17'd59605: data = 8'h0a;
      17'd59606: data = 8'h0a;
      17'd59607: data = 8'h0a;
      17'd59608: data = 8'h0c;
      17'd59609: data = 8'h0c;
      17'd59610: data = 8'h09;
      17'd59611: data = 8'h09;
      17'd59612: data = 8'h0a;
      17'd59613: data = 8'h06;
      17'd59614: data = 8'h01;
      17'd59615: data = 8'h04;
      17'd59616: data = 8'h06;
      17'd59617: data = 8'h0d;
      17'd59618: data = 8'h0d;
      17'd59619: data = 8'h09;
      17'd59620: data = 8'h04;
      17'd59621: data = 8'h02;
      17'd59622: data = 8'h02;
      17'd59623: data = 8'hfd;
      17'd59624: data = 8'hfd;
      17'd59625: data = 8'h00;
      17'd59626: data = 8'h02;
      17'd59627: data = 8'h00;
      17'd59628: data = 8'hfe;
      17'd59629: data = 8'hfe;
      17'd59630: data = 8'h01;
      17'd59631: data = 8'h01;
      17'd59632: data = 8'hfc;
      17'd59633: data = 8'hfe;
      17'd59634: data = 8'h01;
      17'd59635: data = 8'h00;
      17'd59636: data = 8'hfe;
      17'd59637: data = 8'h04;
      17'd59638: data = 8'h05;
      17'd59639: data = 8'h05;
      17'd59640: data = 8'h0a;
      17'd59641: data = 8'h06;
      17'd59642: data = 8'h04;
      17'd59643: data = 8'h05;
      17'd59644: data = 8'h0a;
      17'd59645: data = 8'h09;
      17'd59646: data = 8'h06;
      17'd59647: data = 8'h09;
      17'd59648: data = 8'h09;
      17'd59649: data = 8'h09;
      17'd59650: data = 8'h04;
      17'd59651: data = 8'h01;
      17'd59652: data = 8'h04;
      17'd59653: data = 8'h0a;
      17'd59654: data = 8'h04;
      17'd59655: data = 8'h04;
      17'd59656: data = 8'h0c;
      17'd59657: data = 8'h0c;
      17'd59658: data = 8'h0d;
      17'd59659: data = 8'h0d;
      17'd59660: data = 8'h0d;
      17'd59661: data = 8'h11;
      17'd59662: data = 8'h0c;
      17'd59663: data = 8'h09;
      17'd59664: data = 8'h05;
      17'd59665: data = 8'h04;
      17'd59666: data = 8'h04;
      17'd59667: data = 8'h02;
      17'd59668: data = 8'h01;
      17'd59669: data = 8'hfe;
      17'd59670: data = 8'h00;
      17'd59671: data = 8'hfe;
      17'd59672: data = 8'hfa;
      17'd59673: data = 8'hfa;
      17'd59674: data = 8'hf9;
      17'd59675: data = 8'hf9;
      17'd59676: data = 8'hfa;
      17'd59677: data = 8'hf6;
      17'd59678: data = 8'hf5;
      17'd59679: data = 8'hf6;
      17'd59680: data = 8'hf9;
      17'd59681: data = 8'hf9;
      17'd59682: data = 8'hf9;
      17'd59683: data = 8'hf9;
      17'd59684: data = 8'hf6;
      17'd59685: data = 8'hf5;
      17'd59686: data = 8'hf4;
      17'd59687: data = 8'hf2;
      17'd59688: data = 8'hf5;
      17'd59689: data = 8'hf9;
      17'd59690: data = 8'hfc;
      17'd59691: data = 8'hfa;
      17'd59692: data = 8'hfc;
      17'd59693: data = 8'hfa;
      17'd59694: data = 8'hf9;
      17'd59695: data = 8'hfa;
      17'd59696: data = 8'hf9;
      17'd59697: data = 8'hfa;
      17'd59698: data = 8'hf9;
      17'd59699: data = 8'hf9;
      17'd59700: data = 8'hfc;
      17'd59701: data = 8'hfe;
      17'd59702: data = 8'h00;
      17'd59703: data = 8'hfe;
      17'd59704: data = 8'h00;
      17'd59705: data = 8'h02;
      17'd59706: data = 8'h00;
      17'd59707: data = 8'h04;
      17'd59708: data = 8'h05;
      17'd59709: data = 8'h05;
      17'd59710: data = 8'h0a;
      17'd59711: data = 8'h0c;
      17'd59712: data = 8'h0a;
      17'd59713: data = 8'h09;
      17'd59714: data = 8'h09;
      17'd59715: data = 8'h05;
      17'd59716: data = 8'h06;
      17'd59717: data = 8'h05;
      17'd59718: data = 8'h02;
      17'd59719: data = 8'h01;
      17'd59720: data = 8'h02;
      17'd59721: data = 8'h05;
      17'd59722: data = 8'h04;
      17'd59723: data = 8'h05;
      17'd59724: data = 8'h06;
      17'd59725: data = 8'h04;
      17'd59726: data = 8'h04;
      17'd59727: data = 8'h01;
      17'd59728: data = 8'h00;
      17'd59729: data = 8'h01;
      17'd59730: data = 8'h01;
      17'd59731: data = 8'h01;
      17'd59732: data = 8'h00;
      17'd59733: data = 8'h02;
      17'd59734: data = 8'h05;
      17'd59735: data = 8'h04;
      17'd59736: data = 8'h01;
      17'd59737: data = 8'h02;
      17'd59738: data = 8'h00;
      17'd59739: data = 8'hfe;
      17'd59740: data = 8'hfe;
      17'd59741: data = 8'hfd;
      17'd59742: data = 8'hfe;
      17'd59743: data = 8'hfd;
      17'd59744: data = 8'hfe;
      17'd59745: data = 8'hfd;
      17'd59746: data = 8'hfc;
      17'd59747: data = 8'hfc;
      17'd59748: data = 8'hfa;
      17'd59749: data = 8'hfa;
      17'd59750: data = 8'hfa;
      17'd59751: data = 8'hf6;
      17'd59752: data = 8'hfd;
      17'd59753: data = 8'hfd;
      17'd59754: data = 8'hfa;
      17'd59755: data = 8'hfa;
      17'd59756: data = 8'hfc;
      17'd59757: data = 8'hfe;
      17'd59758: data = 8'hfa;
      17'd59759: data = 8'hfa;
      17'd59760: data = 8'hf9;
      17'd59761: data = 8'hf9;
      17'd59762: data = 8'hf9;
      17'd59763: data = 8'hf4;
      17'd59764: data = 8'hf5;
      17'd59765: data = 8'hf6;
      17'd59766: data = 8'hf5;
      17'd59767: data = 8'hf4;
      17'd59768: data = 8'hf4;
      17'd59769: data = 8'hf4;
      17'd59770: data = 8'hf1;
      17'd59771: data = 8'hf1;
      17'd59772: data = 8'hf2;
      17'd59773: data = 8'hf1;
      17'd59774: data = 8'hef;
      17'd59775: data = 8'hef;
      17'd59776: data = 8'hef;
      17'd59777: data = 8'hed;
      17'd59778: data = 8'hed;
      17'd59779: data = 8'hec;
      17'd59780: data = 8'hed;
      17'd59781: data = 8'hef;
      17'd59782: data = 8'hef;
      17'd59783: data = 8'hef;
      17'd59784: data = 8'hf1;
      17'd59785: data = 8'hf4;
      17'd59786: data = 8'hf2;
      17'd59787: data = 8'hf2;
      17'd59788: data = 8'hf1;
      17'd59789: data = 8'hed;
      17'd59790: data = 8'hed;
      17'd59791: data = 8'hed;
      17'd59792: data = 8'hed;
      17'd59793: data = 8'hef;
      17'd59794: data = 8'hef;
      17'd59795: data = 8'hef;
      17'd59796: data = 8'hf1;
      17'd59797: data = 8'hf2;
      17'd59798: data = 8'hf2;
      17'd59799: data = 8'hf4;
      17'd59800: data = 8'hf4;
      17'd59801: data = 8'hf6;
      17'd59802: data = 8'hf9;
      17'd59803: data = 8'hf5;
      17'd59804: data = 8'hf9;
      17'd59805: data = 8'hfc;
      17'd59806: data = 8'hfd;
      17'd59807: data = 8'hfe;
      17'd59808: data = 8'h00;
      17'd59809: data = 8'h01;
      17'd59810: data = 8'h01;
      17'd59811: data = 8'h02;
      17'd59812: data = 8'h04;
      17'd59813: data = 8'h05;
      17'd59814: data = 8'h05;
      17'd59815: data = 8'h09;
      17'd59816: data = 8'h0c;
      17'd59817: data = 8'h0a;
      17'd59818: data = 8'h0c;
      17'd59819: data = 8'h0d;
      17'd59820: data = 8'h0d;
      17'd59821: data = 8'h0e;
      17'd59822: data = 8'h0d;
      17'd59823: data = 8'h0a;
      17'd59824: data = 8'h0d;
      17'd59825: data = 8'h0e;
      17'd59826: data = 8'h0d;
      17'd59827: data = 8'h11;
      17'd59828: data = 8'h11;
      17'd59829: data = 8'h12;
      17'd59830: data = 8'h11;
      17'd59831: data = 8'h11;
      17'd59832: data = 8'h12;
      17'd59833: data = 8'h0e;
      17'd59834: data = 8'h0e;
      17'd59835: data = 8'h11;
      17'd59836: data = 8'h0e;
      17'd59837: data = 8'h11;
      17'd59838: data = 8'h0c;
      17'd59839: data = 8'h04;
      17'd59840: data = 8'h04;
      17'd59841: data = 8'h09;
      17'd59842: data = 8'h0c;
      17'd59843: data = 8'h09;
      17'd59844: data = 8'h04;
      17'd59845: data = 8'h06;
      17'd59846: data = 8'h0e;
      17'd59847: data = 8'h11;
      17'd59848: data = 8'h0a;
      17'd59849: data = 8'h04;
      17'd59850: data = 8'h06;
      17'd59851: data = 8'h0c;
      17'd59852: data = 8'h0c;
      17'd59853: data = 8'h01;
      17'd59854: data = 8'hfc;
      17'd59855: data = 8'h01;
      17'd59856: data = 8'h09;
      17'd59857: data = 8'h06;
      17'd59858: data = 8'h01;
      17'd59859: data = 8'hfd;
      17'd59860: data = 8'hfd;
      17'd59861: data = 8'h02;
      17'd59862: data = 8'h04;
      17'd59863: data = 8'h02;
      17'd59864: data = 8'h00;
      17'd59865: data = 8'h00;
      17'd59866: data = 8'h04;
      17'd59867: data = 8'h04;
      17'd59868: data = 8'h02;
      17'd59869: data = 8'h00;
      17'd59870: data = 8'h01;
      17'd59871: data = 8'h02;
      17'd59872: data = 8'h02;
      17'd59873: data = 8'h00;
      17'd59874: data = 8'hfd;
      17'd59875: data = 8'hfc;
      17'd59876: data = 8'hfd;
      17'd59877: data = 8'hfe;
      17'd59878: data = 8'hfd;
      17'd59879: data = 8'h01;
      17'd59880: data = 8'h02;
      17'd59881: data = 8'h04;
      17'd59882: data = 8'h04;
      17'd59883: data = 8'h01;
      17'd59884: data = 8'h02;
      17'd59885: data = 8'h01;
      17'd59886: data = 8'hfe;
      17'd59887: data = 8'hfd;
      17'd59888: data = 8'h01;
      17'd59889: data = 8'h04;
      17'd59890: data = 8'h04;
      17'd59891: data = 8'h01;
      17'd59892: data = 8'h04;
      17'd59893: data = 8'h09;
      17'd59894: data = 8'h06;
      17'd59895: data = 8'h05;
      17'd59896: data = 8'h05;
      17'd59897: data = 8'h09;
      17'd59898: data = 8'h05;
      17'd59899: data = 8'h05;
      17'd59900: data = 8'h09;
      17'd59901: data = 8'h0a;
      17'd59902: data = 8'h0a;
      17'd59903: data = 8'h0a;
      17'd59904: data = 8'h0c;
      17'd59905: data = 8'h09;
      17'd59906: data = 8'h05;
      17'd59907: data = 8'h05;
      17'd59908: data = 8'h06;
      17'd59909: data = 8'h05;
      17'd59910: data = 8'h04;
      17'd59911: data = 8'h05;
      17'd59912: data = 8'h09;
      17'd59913: data = 8'h04;
      17'd59914: data = 8'h04;
      17'd59915: data = 8'h09;
      17'd59916: data = 8'h0a;
      17'd59917: data = 8'h02;
      17'd59918: data = 8'hfe;
      17'd59919: data = 8'hfe;
      17'd59920: data = 8'hfd;
      17'd59921: data = 8'hfc;
      17'd59922: data = 8'hf9;
      17'd59923: data = 8'hfc;
      17'd59924: data = 8'hfd;
      17'd59925: data = 8'hfc;
      17'd59926: data = 8'hfd;
      17'd59927: data = 8'hfa;
      17'd59928: data = 8'hf6;
      17'd59929: data = 8'hf5;
      17'd59930: data = 8'hf4;
      17'd59931: data = 8'hf2;
      17'd59932: data = 8'hf5;
      17'd59933: data = 8'hf4;
      17'd59934: data = 8'hf4;
      17'd59935: data = 8'hf5;
      17'd59936: data = 8'hf4;
      17'd59937: data = 8'hf4;
      17'd59938: data = 8'hf4;
      17'd59939: data = 8'hf4;
      17'd59940: data = 8'hf2;
      17'd59941: data = 8'hef;
      17'd59942: data = 8'hf4;
      17'd59943: data = 8'hf6;
      17'd59944: data = 8'hf6;
      17'd59945: data = 8'hf9;
      17'd59946: data = 8'hf9;
      17'd59947: data = 8'hf9;
      17'd59948: data = 8'hf6;
      17'd59949: data = 8'hf6;
      17'd59950: data = 8'hf9;
      17'd59951: data = 8'hf9;
      17'd59952: data = 8'hfd;
      17'd59953: data = 8'hfe;
      17'd59954: data = 8'h00;
      17'd59955: data = 8'h01;
      17'd59956: data = 8'h01;
      17'd59957: data = 8'h01;
      17'd59958: data = 8'h01;
      17'd59959: data = 8'h00;
      17'd59960: data = 8'hfe;
      17'd59961: data = 8'hfd;
      17'd59962: data = 8'hfd;
      17'd59963: data = 8'h00;
      17'd59964: data = 8'h01;
      17'd59965: data = 8'h02;
      17'd59966: data = 8'h02;
      17'd59967: data = 8'h04;
      17'd59968: data = 8'h02;
      17'd59969: data = 8'h04;
      17'd59970: data = 8'h02;
      17'd59971: data = 8'h00;
      17'd59972: data = 8'h00;
      17'd59973: data = 8'h00;
      17'd59974: data = 8'h01;
      17'd59975: data = 8'h01;
      17'd59976: data = 8'h00;
      17'd59977: data = 8'h00;
      17'd59978: data = 8'h00;
      17'd59979: data = 8'h00;
      17'd59980: data = 8'hfe;
      17'd59981: data = 8'hfe;
      17'd59982: data = 8'hfd;
      17'd59983: data = 8'hfe;
      17'd59984: data = 8'h00;
      17'd59985: data = 8'hfe;
      17'd59986: data = 8'hfe;
      17'd59987: data = 8'h00;
      17'd59988: data = 8'h01;
      17'd59989: data = 8'hfe;
      17'd59990: data = 8'hfe;
      17'd59991: data = 8'hfe;
      17'd59992: data = 8'hfc;
      17'd59993: data = 8'hfc;
      17'd59994: data = 8'hfa;
      17'd59995: data = 8'hf9;
      17'd59996: data = 8'hfc;
      17'd59997: data = 8'hfa;
      17'd59998: data = 8'hfc;
      17'd59999: data = 8'hfc;
      17'd60000: data = 8'hfa;
      17'd60001: data = 8'hfc;
      17'd60002: data = 8'hfe;
      17'd60003: data = 8'hfd;
      17'd60004: data = 8'hfe;
      17'd60005: data = 8'hfc;
      17'd60006: data = 8'hf9;
      17'd60007: data = 8'hfa;
      17'd60008: data = 8'hf6;
      17'd60009: data = 8'hf6;
      17'd60010: data = 8'hf4;
      17'd60011: data = 8'hf5;
      17'd60012: data = 8'hf5;
      17'd60013: data = 8'hf2;
      17'd60014: data = 8'hf4;
      17'd60015: data = 8'hf5;
      17'd60016: data = 8'hf2;
      17'd60017: data = 8'hf4;
      17'd60018: data = 8'hf5;
      17'd60019: data = 8'hf1;
      17'd60020: data = 8'hf1;
      17'd60021: data = 8'hef;
      17'd60022: data = 8'hec;
      17'd60023: data = 8'heb;
      17'd60024: data = 8'hed;
      17'd60025: data = 8'heb;
      17'd60026: data = 8'heb;
      17'd60027: data = 8'hec;
      17'd60028: data = 8'hec;
      17'd60029: data = 8'hef;
      17'd60030: data = 8'hf1;
      17'd60031: data = 8'hef;
      17'd60032: data = 8'hec;
      17'd60033: data = 8'hec;
      17'd60034: data = 8'hed;
      17'd60035: data = 8'hef;
      17'd60036: data = 8'hef;
      17'd60037: data = 8'hf1;
      17'd60038: data = 8'hf4;
      17'd60039: data = 8'hf4;
      17'd60040: data = 8'hf4;
      17'd60041: data = 8'hf1;
      17'd60042: data = 8'hf1;
      17'd60043: data = 8'hf2;
      17'd60044: data = 8'hf2;
      17'd60045: data = 8'hf5;
      17'd60046: data = 8'hf9;
      17'd60047: data = 8'hfa;
      17'd60048: data = 8'hfd;
      17'd60049: data = 8'hfd;
      17'd60050: data = 8'hfd;
      17'd60051: data = 8'hfe;
      17'd60052: data = 8'h00;
      17'd60053: data = 8'h00;
      17'd60054: data = 8'h01;
      17'd60055: data = 8'h01;
      17'd60056: data = 8'h01;
      17'd60057: data = 8'h02;
      17'd60058: data = 8'h05;
      17'd60059: data = 8'h05;
      17'd60060: data = 8'h05;
      17'd60061: data = 8'h05;
      17'd60062: data = 8'h05;
      17'd60063: data = 8'h06;
      17'd60064: data = 8'h09;
      17'd60065: data = 8'h06;
      17'd60066: data = 8'h06;
      17'd60067: data = 8'h0d;
      17'd60068: data = 8'h0e;
      17'd60069: data = 8'h0a;
      17'd60070: data = 8'h0d;
      17'd60071: data = 8'h12;
      17'd60072: data = 8'h12;
      17'd60073: data = 8'h11;
      17'd60074: data = 8'h09;
      17'd60075: data = 8'h06;
      17'd60076: data = 8'h0c;
      17'd60077: data = 8'h0d;
      17'd60078: data = 8'h09;
      17'd60079: data = 8'h06;
      17'd60080: data = 8'h0c;
      17'd60081: data = 8'h12;
      17'd60082: data = 8'h11;
      17'd60083: data = 8'h0c;
      17'd60084: data = 8'h09;
      17'd60085: data = 8'h0a;
      17'd60086: data = 8'h0e;
      17'd60087: data = 8'h11;
      17'd60088: data = 8'h0c;
      17'd60089: data = 8'h06;
      17'd60090: data = 8'h0c;
      17'd60091: data = 8'h0d;
      17'd60092: data = 8'h0a;
      17'd60093: data = 8'h09;
      17'd60094: data = 8'h09;
      17'd60095: data = 8'h09;
      17'd60096: data = 8'h0a;
      17'd60097: data = 8'h0c;
      17'd60098: data = 8'h09;
      17'd60099: data = 8'h09;
      17'd60100: data = 8'h09;
      17'd60101: data = 8'h06;
      17'd60102: data = 8'h0c;
      17'd60103: data = 8'h0e;
      17'd60104: data = 8'h09;
      17'd60105: data = 8'h04;
      17'd60106: data = 8'h01;
      17'd60107: data = 8'h04;
      17'd60108: data = 8'h06;
      17'd60109: data = 8'h04;
      17'd60110: data = 8'hfd;
      17'd60111: data = 8'h01;
      17'd60112: data = 8'h09;
      17'd60113: data = 8'h05;
      17'd60114: data = 8'h01;
      17'd60115: data = 8'h00;
      17'd60116: data = 8'h04;
      17'd60117: data = 8'h05;
      17'd60118: data = 8'h04;
      17'd60119: data = 8'h02;
      17'd60120: data = 8'h00;
      17'd60121: data = 8'h00;
      17'd60122: data = 8'h02;
      17'd60123: data = 8'h05;
      17'd60124: data = 8'h05;
      17'd60125: data = 8'h02;
      17'd60126: data = 8'h01;
      17'd60127: data = 8'h00;
      17'd60128: data = 8'hfd;
      17'd60129: data = 8'hfe;
      17'd60130: data = 8'h01;
      17'd60131: data = 8'hfe;
      17'd60132: data = 8'hfd;
      17'd60133: data = 8'hfe;
      17'd60134: data = 8'h02;
      17'd60135: data = 8'h01;
      17'd60136: data = 8'hfd;
      17'd60137: data = 8'hfe;
      17'd60138: data = 8'h01;
      17'd60139: data = 8'h00;
      17'd60140: data = 8'hfd;
      17'd60141: data = 8'hfd;
      17'd60142: data = 8'h01;
      17'd60143: data = 8'h02;
      17'd60144: data = 8'h04;
      17'd60145: data = 8'h04;
      17'd60146: data = 8'h04;
      17'd60147: data = 8'h01;
      17'd60148: data = 8'h00;
      17'd60149: data = 8'h01;
      17'd60150: data = 8'h02;
      17'd60151: data = 8'h06;
      17'd60152: data = 8'h09;
      17'd60153: data = 8'h09;
      17'd60154: data = 8'h09;
      17'd60155: data = 8'h09;
      17'd60156: data = 8'h09;
      17'd60157: data = 8'h05;
      17'd60158: data = 8'h05;
      17'd60159: data = 8'h04;
      17'd60160: data = 8'h05;
      17'd60161: data = 8'h06;
      17'd60162: data = 8'h06;
      17'd60163: data = 8'h09;
      17'd60164: data = 8'h0c;
      17'd60165: data = 8'h0c;
      17'd60166: data = 8'h0c;
      17'd60167: data = 8'h0c;
      17'd60168: data = 8'h0c;
      17'd60169: data = 8'h0c;
      17'd60170: data = 8'h0c;
      17'd60171: data = 8'h0a;
      17'd60172: data = 8'h0a;
      17'd60173: data = 8'h0c;
      17'd60174: data = 8'h0a;
      17'd60175: data = 8'h0a;
      17'd60176: data = 8'h06;
      17'd60177: data = 8'h06;
      17'd60178: data = 8'h04;
      17'd60179: data = 8'h00;
      17'd60180: data = 8'hfe;
      17'd60181: data = 8'hfd;
      17'd60182: data = 8'hfd;
      17'd60183: data = 8'hfe;
      17'd60184: data = 8'hfd;
      17'd60185: data = 8'h00;
      17'd60186: data = 8'hfe;
      17'd60187: data = 8'hfc;
      17'd60188: data = 8'hfa;
      17'd60189: data = 8'hf6;
      17'd60190: data = 8'hf5;
      17'd60191: data = 8'hf2;
      17'd60192: data = 8'hf2;
      17'd60193: data = 8'hf1;
      17'd60194: data = 8'hf1;
      17'd60195: data = 8'hf5;
      17'd60196: data = 8'hf6;
      17'd60197: data = 8'hf6;
      17'd60198: data = 8'hf5;
      17'd60199: data = 8'hf4;
      17'd60200: data = 8'hf4;
      17'd60201: data = 8'hf1;
      17'd60202: data = 8'hed;
      17'd60203: data = 8'hec;
      17'd60204: data = 8'hef;
      17'd60205: data = 8'hf1;
      17'd60206: data = 8'hf2;
      17'd60207: data = 8'hf2;
      17'd60208: data = 8'hf2;
      17'd60209: data = 8'hf2;
      17'd60210: data = 8'hf1;
      17'd60211: data = 8'hf1;
      17'd60212: data = 8'hf2;
      17'd60213: data = 8'hf2;
      17'd60214: data = 8'hf4;
      17'd60215: data = 8'hf6;
      17'd60216: data = 8'hf6;
      17'd60217: data = 8'hf6;
      17'd60218: data = 8'hf9;
      17'd60219: data = 8'hfc;
      17'd60220: data = 8'hfa;
      17'd60221: data = 8'hf6;
      17'd60222: data = 8'hf9;
      17'd60223: data = 8'hf6;
      17'd60224: data = 8'hf5;
      17'd60225: data = 8'hf6;
      17'd60226: data = 8'hf9;
      17'd60227: data = 8'hfa;
      17'd60228: data = 8'hfa;
      17'd60229: data = 8'hfa;
      17'd60230: data = 8'hfd;
      17'd60231: data = 8'hfc;
      17'd60232: data = 8'hfa;
      17'd60233: data = 8'hfc;
      17'd60234: data = 8'hfd;
      17'd60235: data = 8'hfe;
      17'd60236: data = 8'hfe;
      17'd60237: data = 8'h00;
      17'd60238: data = 8'h00;
      17'd60239: data = 8'hfe;
      17'd60240: data = 8'hfd;
      17'd60241: data = 8'hfd;
      17'd60242: data = 8'hfd;
      17'd60243: data = 8'hfc;
      17'd60244: data = 8'hfc;
      17'd60245: data = 8'hfd;
      17'd60246: data = 8'hfd;
      17'd60247: data = 8'hfe;
      17'd60248: data = 8'h01;
      17'd60249: data = 8'h02;
      17'd60250: data = 8'h02;
      17'd60251: data = 8'h00;
      17'd60252: data = 8'h00;
      17'd60253: data = 8'h00;
      17'd60254: data = 8'hfd;
      17'd60255: data = 8'hfc;
      17'd60256: data = 8'hfc;
      17'd60257: data = 8'hfd;
      17'd60258: data = 8'hfe;
      17'd60259: data = 8'hfd;
      17'd60260: data = 8'hfe;
      17'd60261: data = 8'hfe;
      17'd60262: data = 8'hfe;
      17'd60263: data = 8'hfe;
      17'd60264: data = 8'hfd;
      17'd60265: data = 8'hfe;
      17'd60266: data = 8'hfe;
      17'd60267: data = 8'hfe;
      17'd60268: data = 8'h00;
      17'd60269: data = 8'h00;
      17'd60270: data = 8'hfe;
      17'd60271: data = 8'hfd;
      17'd60272: data = 8'hfd;
      17'd60273: data = 8'hfc;
      17'd60274: data = 8'hfc;
      17'd60275: data = 8'hfc;
      17'd60276: data = 8'hfa;
      17'd60277: data = 8'hfc;
      17'd60278: data = 8'hfd;
      17'd60279: data = 8'hfd;
      17'd60280: data = 8'h00;
      17'd60281: data = 8'hfe;
      17'd60282: data = 8'hfd;
      17'd60283: data = 8'hfc;
      17'd60284: data = 8'hfc;
      17'd60285: data = 8'hfc;
      17'd60286: data = 8'hfc;
      17'd60287: data = 8'hfa;
      17'd60288: data = 8'hfa;
      17'd60289: data = 8'hfc;
      17'd60290: data = 8'hfc;
      17'd60291: data = 8'hfc;
      17'd60292: data = 8'hfc;
      17'd60293: data = 8'hfc;
      17'd60294: data = 8'hfa;
      17'd60295: data = 8'hfa;
      17'd60296: data = 8'hfa;
      17'd60297: data = 8'hfa;
      17'd60298: data = 8'hf6;
      17'd60299: data = 8'hf6;
      17'd60300: data = 8'hf9;
      17'd60301: data = 8'hfa;
      17'd60302: data = 8'hf9;
      17'd60303: data = 8'hf9;
      17'd60304: data = 8'hf9;
      17'd60305: data = 8'hf9;
      17'd60306: data = 8'hf6;
      17'd60307: data = 8'hf9;
      17'd60308: data = 8'hf6;
      17'd60309: data = 8'hf6;
      17'd60310: data = 8'hfa;
      17'd60311: data = 8'hf9;
      17'd60312: data = 8'hf6;
      17'd60313: data = 8'hf6;
      17'd60314: data = 8'hfa;
      17'd60315: data = 8'hfc;
      17'd60316: data = 8'hfa;
      17'd60317: data = 8'hfc;
      17'd60318: data = 8'hfd;
      17'd60319: data = 8'hfd;
      17'd60320: data = 8'hfd;
      17'd60321: data = 8'hfd;
      17'd60322: data = 8'h01;
      17'd60323: data = 8'h04;
      17'd60324: data = 8'h01;
      17'd60325: data = 8'hfe;
      17'd60326: data = 8'hfe;
      17'd60327: data = 8'hfe;
      17'd60328: data = 8'h00;
      17'd60329: data = 8'h02;
      17'd60330: data = 8'h01;
      17'd60331: data = 8'h02;
      17'd60332: data = 8'h05;
      17'd60333: data = 8'h05;
      17'd60334: data = 8'h05;
      17'd60335: data = 8'h02;
      17'd60336: data = 8'h04;
      17'd60337: data = 8'h0a;
      17'd60338: data = 8'h0a;
      17'd60339: data = 8'h09;
      17'd60340: data = 8'h0c;
      17'd60341: data = 8'h0d;
      17'd60342: data = 8'h0d;
      17'd60343: data = 8'h11;
      17'd60344: data = 8'h13;
      17'd60345: data = 8'h0d;
      17'd60346: data = 8'h0c;
      17'd60347: data = 8'h0d;
      17'd60348: data = 8'h0d;
      17'd60349: data = 8'h0c;
      17'd60350: data = 8'h0c;
      17'd60351: data = 8'h0c;
      17'd60352: data = 8'h0e;
      17'd60353: data = 8'h0e;
      17'd60354: data = 8'h0d;
      17'd60355: data = 8'h0d;
      17'd60356: data = 8'h0c;
      17'd60357: data = 8'h0c;
      17'd60358: data = 8'h0d;
      17'd60359: data = 8'h0c;
      17'd60360: data = 8'h0c;
      17'd60361: data = 8'h0c;
      17'd60362: data = 8'h0d;
      17'd60363: data = 8'h0c;
      17'd60364: data = 8'h0a;
      17'd60365: data = 8'h0d;
      17'd60366: data = 8'h0d;
      17'd60367: data = 8'h0a;
      17'd60368: data = 8'h0d;
      17'd60369: data = 8'h09;
      17'd60370: data = 8'h06;
      17'd60371: data = 8'h06;
      17'd60372: data = 8'h06;
      17'd60373: data = 8'h06;
      17'd60374: data = 8'h05;
      17'd60375: data = 8'h05;
      17'd60376: data = 8'h02;
      17'd60377: data = 8'h04;
      17'd60378: data = 8'h05;
      17'd60379: data = 8'h04;
      17'd60380: data = 8'h04;
      17'd60381: data = 8'h02;
      17'd60382: data = 8'h02;
      17'd60383: data = 8'h04;
      17'd60384: data = 8'h02;
      17'd60385: data = 8'h04;
      17'd60386: data = 8'h05;
      17'd60387: data = 8'h05;
      17'd60388: data = 8'h06;
      17'd60389: data = 8'h05;
      17'd60390: data = 8'h05;
      17'd60391: data = 8'h04;
      17'd60392: data = 8'h06;
      17'd60393: data = 8'h04;
      17'd60394: data = 8'h02;
      17'd60395: data = 8'h02;
      17'd60396: data = 8'h01;
      17'd60397: data = 8'h00;
      17'd60398: data = 8'h01;
      17'd60399: data = 8'h00;
      17'd60400: data = 8'h00;
      17'd60401: data = 8'h01;
      17'd60402: data = 8'h02;
      17'd60403: data = 8'h02;
      17'd60404: data = 8'h01;
      17'd60405: data = 8'h01;
      17'd60406: data = 8'h01;
      17'd60407: data = 8'h01;
      17'd60408: data = 8'h00;
      17'd60409: data = 8'hfe;
      17'd60410: data = 8'hfc;
      17'd60411: data = 8'hfd;
      17'd60412: data = 8'h02;
      17'd60413: data = 8'h02;
      17'd60414: data = 8'h02;
      17'd60415: data = 8'h02;
      17'd60416: data = 8'h01;
      17'd60417: data = 8'h02;
      17'd60418: data = 8'h00;
      17'd60419: data = 8'hfd;
      17'd60420: data = 8'hfd;
      17'd60421: data = 8'hfe;
      17'd60422: data = 8'hfd;
      17'd60423: data = 8'hfd;
      17'd60424: data = 8'hfc;
      17'd60425: data = 8'hfc;
      17'd60426: data = 8'hfd;
      17'd60427: data = 8'hfc;
      17'd60428: data = 8'hfa;
      17'd60429: data = 8'hfc;
      17'd60430: data = 8'hfc;
      17'd60431: data = 8'hfc;
      17'd60432: data = 8'hfe;
      17'd60433: data = 8'hfe;
      17'd60434: data = 8'h00;
      17'd60435: data = 8'hfe;
      17'd60436: data = 8'h00;
      17'd60437: data = 8'hfe;
      17'd60438: data = 8'hfd;
      17'd60439: data = 8'hfc;
      17'd60440: data = 8'hfa;
      17'd60441: data = 8'hfc;
      17'd60442: data = 8'hfa;
      17'd60443: data = 8'hfc;
      17'd60444: data = 8'hfa;
      17'd60445: data = 8'hf9;
      17'd60446: data = 8'hfa;
      17'd60447: data = 8'hfd;
      17'd60448: data = 8'hf9;
      17'd60449: data = 8'hf9;
      17'd60450: data = 8'hfa;
      17'd60451: data = 8'hfa;
      17'd60452: data = 8'hf9;
      17'd60453: data = 8'hfc;
      17'd60454: data = 8'hfc;
      17'd60455: data = 8'hf9;
      17'd60456: data = 8'hf6;
      17'd60457: data = 8'hf6;
      17'd60458: data = 8'hf9;
      17'd60459: data = 8'hf5;
      17'd60460: data = 8'hf6;
      17'd60461: data = 8'hf6;
      17'd60462: data = 8'hf9;
      17'd60463: data = 8'hf9;
      17'd60464: data = 8'hfc;
      17'd60465: data = 8'hfa;
      17'd60466: data = 8'hf9;
      17'd60467: data = 8'hf9;
      17'd60468: data = 8'hf9;
      17'd60469: data = 8'hf9;
      17'd60470: data = 8'hf6;
      17'd60471: data = 8'hf9;
      17'd60472: data = 8'hfa;
      17'd60473: data = 8'hf6;
      17'd60474: data = 8'hf9;
      17'd60475: data = 8'hf9;
      17'd60476: data = 8'hf6;
      17'd60477: data = 8'hf9;
      17'd60478: data = 8'hf9;
      17'd60479: data = 8'hf6;
      17'd60480: data = 8'hf5;
      17'd60481: data = 8'hf6;
      17'd60482: data = 8'hf5;
      17'd60483: data = 8'hf4;
      17'd60484: data = 8'hf4;
      17'd60485: data = 8'hf6;
      17'd60486: data = 8'hf6;
      17'd60487: data = 8'hf5;
      17'd60488: data = 8'hf4;
      17'd60489: data = 8'hf2;
      17'd60490: data = 8'hf4;
      17'd60491: data = 8'hf4;
      17'd60492: data = 8'hf4;
      17'd60493: data = 8'hf5;
      17'd60494: data = 8'hf2;
      17'd60495: data = 8'hf4;
      17'd60496: data = 8'hf4;
      17'd60497: data = 8'hf4;
      17'd60498: data = 8'hf4;
      17'd60499: data = 8'hf4;
      17'd60500: data = 8'hf4;
      17'd60501: data = 8'hf2;
      17'd60502: data = 8'hf5;
      17'd60503: data = 8'hf4;
      17'd60504: data = 8'hf2;
      17'd60505: data = 8'hf1;
      17'd60506: data = 8'hf1;
      17'd60507: data = 8'hf4;
      17'd60508: data = 8'hf9;
      17'd60509: data = 8'hf9;
      17'd60510: data = 8'hf9;
      17'd60511: data = 8'hf9;
      17'd60512: data = 8'hf9;
      17'd60513: data = 8'hf9;
      17'd60514: data = 8'hf9;
      17'd60515: data = 8'hfa;
      17'd60516: data = 8'hfa;
      17'd60517: data = 8'hfa;
      17'd60518: data = 8'hfa;
      17'd60519: data = 8'hf9;
      17'd60520: data = 8'hfd;
      17'd60521: data = 8'hfd;
      17'd60522: data = 8'hfd;
      17'd60523: data = 8'h00;
      17'd60524: data = 8'h01;
      17'd60525: data = 8'h00;
      17'd60526: data = 8'h02;
      17'd60527: data = 8'h02;
      17'd60528: data = 8'h01;
      17'd60529: data = 8'h02;
      17'd60530: data = 8'h04;
      17'd60531: data = 8'h05;
      17'd60532: data = 8'h02;
      17'd60533: data = 8'h02;
      17'd60534: data = 8'h02;
      17'd60535: data = 8'h04;
      17'd60536: data = 8'h06;
      17'd60537: data = 8'h04;
      17'd60538: data = 8'h05;
      17'd60539: data = 8'h06;
      17'd60540: data = 8'h05;
      17'd60541: data = 8'h05;
      17'd60542: data = 8'h06;
      17'd60543: data = 8'h05;
      17'd60544: data = 8'h06;
      17'd60545: data = 8'h05;
      17'd60546: data = 8'h05;
      17'd60547: data = 8'h05;
      17'd60548: data = 8'h02;
      17'd60549: data = 8'h02;
      17'd60550: data = 8'h05;
      17'd60551: data = 8'h02;
      17'd60552: data = 8'h01;
      17'd60553: data = 8'h02;
      17'd60554: data = 8'h02;
      17'd60555: data = 8'h05;
      17'd60556: data = 8'h01;
      17'd60557: data = 8'h04;
      17'd60558: data = 8'h06;
      17'd60559: data = 8'h05;
      17'd60560: data = 8'h02;
      17'd60561: data = 8'h04;
      17'd60562: data = 8'h02;
      17'd60563: data = 8'h02;
      17'd60564: data = 8'h05;
      17'd60565: data = 8'h01;
      17'd60566: data = 8'h01;
      17'd60567: data = 8'h01;
      17'd60568: data = 8'h02;
      17'd60569: data = 8'h01;
      17'd60570: data = 8'h01;
      17'd60571: data = 8'h01;
      17'd60572: data = 8'h01;
      17'd60573: data = 8'h01;
      17'd60574: data = 8'h02;
      17'd60575: data = 8'h00;
      17'd60576: data = 8'hfd;
      17'd60577: data = 8'h01;
      17'd60578: data = 8'h02;
      17'd60579: data = 8'h02;
      17'd60580: data = 8'h00;
      17'd60581: data = 8'hfe;
      17'd60582: data = 8'h00;
      17'd60583: data = 8'h00;
      17'd60584: data = 8'h00;
      17'd60585: data = 8'h00;
      17'd60586: data = 8'hfe;
      17'd60587: data = 8'hfe;
      17'd60588: data = 8'h01;
      17'd60589: data = 8'hfe;
      17'd60590: data = 8'hfc;
      17'd60591: data = 8'hfe;
      17'd60592: data = 8'h00;
      17'd60593: data = 8'h01;
      17'd60594: data = 8'hfe;
      17'd60595: data = 8'h00;
      17'd60596: data = 8'hfe;
      17'd60597: data = 8'h00;
      17'd60598: data = 8'h00;
      17'd60599: data = 8'hfe;
      17'd60600: data = 8'h01;
      17'd60601: data = 8'h04;
      17'd60602: data = 8'h02;
      17'd60603: data = 8'h01;
      17'd60604: data = 8'hfd;
      17'd60605: data = 8'hfe;
      17'd60606: data = 8'h01;
      17'd60607: data = 8'hfd;
      17'd60608: data = 8'hfe;
      17'd60609: data = 8'hfe;
      17'd60610: data = 8'hfe;
      17'd60611: data = 8'h01;
      17'd60612: data = 8'h04;
      17'd60613: data = 8'h04;
      17'd60614: data = 8'h04;
      17'd60615: data = 8'h05;
      17'd60616: data = 8'h05;
      17'd60617: data = 8'h01;
      17'd60618: data = 8'h01;
      17'd60619: data = 8'h04;
      17'd60620: data = 8'h02;
      17'd60621: data = 8'h01;
      17'd60622: data = 8'h02;
      17'd60623: data = 8'h01;
      17'd60624: data = 8'h00;
      17'd60625: data = 8'h01;
      17'd60626: data = 8'h01;
      17'd60627: data = 8'h04;
      17'd60628: data = 8'h05;
      17'd60629: data = 8'h0a;
      17'd60630: data = 8'h0c;
      17'd60631: data = 8'h0a;
      17'd60632: data = 8'h0e;
      17'd60633: data = 8'h0c;
      17'd60634: data = 8'h09;
      17'd60635: data = 8'h0d;
      17'd60636: data = 8'h0a;
      17'd60637: data = 8'h06;
      17'd60638: data = 8'h09;
      17'd60639: data = 8'h09;
      17'd60640: data = 8'h0c;
      17'd60641: data = 8'h0e;
      17'd60642: data = 8'h0e;
      17'd60643: data = 8'h0d;
      17'd60644: data = 8'h0e;
      17'd60645: data = 8'h0d;
      17'd60646: data = 8'h0e;
      17'd60647: data = 8'h11;
      17'd60648: data = 8'h0a;
      17'd60649: data = 8'h0e;
      17'd60650: data = 8'h12;
      17'd60651: data = 8'h0c;
      17'd60652: data = 8'h0c;
      17'd60653: data = 8'h0d;
      17'd60654: data = 8'h0a;
      17'd60655: data = 8'h0d;
      17'd60656: data = 8'h0d;
      17'd60657: data = 8'h0c;
      17'd60658: data = 8'h0d;
      17'd60659: data = 8'h0d;
      17'd60660: data = 8'h0c;
      17'd60661: data = 8'h06;
      17'd60662: data = 8'h0a;
      17'd60663: data = 8'h06;
      17'd60664: data = 8'h05;
      17'd60665: data = 8'h05;
      17'd60666: data = 8'h02;
      17'd60667: data = 8'h01;
      17'd60668: data = 8'h00;
      17'd60669: data = 8'hfe;
      17'd60670: data = 8'hfd;
      17'd60671: data = 8'hfd;
      17'd60672: data = 8'hfe;
      17'd60673: data = 8'h01;
      17'd60674: data = 8'hfe;
      17'd60675: data = 8'hfd;
      17'd60676: data = 8'h00;
      17'd60677: data = 8'h01;
      17'd60678: data = 8'h00;
      17'd60679: data = 8'hfc;
      17'd60680: data = 8'hfa;
      17'd60681: data = 8'hfc;
      17'd60682: data = 8'hfa;
      17'd60683: data = 8'hf6;
      17'd60684: data = 8'hf4;
      17'd60685: data = 8'hf5;
      17'd60686: data = 8'hf6;
      17'd60687: data = 8'hf9;
      17'd60688: data = 8'hf9;
      17'd60689: data = 8'hfc;
      17'd60690: data = 8'hfc;
      17'd60691: data = 8'hfa;
      17'd60692: data = 8'hfd;
      17'd60693: data = 8'hfc;
      17'd60694: data = 8'hfa;
      17'd60695: data = 8'hf5;
      17'd60696: data = 8'hf6;
      17'd60697: data = 8'hf9;
      17'd60698: data = 8'hf5;
      17'd60699: data = 8'hf4;
      17'd60700: data = 8'hf2;
      17'd60701: data = 8'hf5;
      17'd60702: data = 8'hf6;
      17'd60703: data = 8'hf9;
      17'd60704: data = 8'hf9;
      17'd60705: data = 8'hf6;
      17'd60706: data = 8'hfa;
      17'd60707: data = 8'hfc;
      17'd60708: data = 8'hfc;
      17'd60709: data = 8'hf9;
      17'd60710: data = 8'hf9;
      17'd60711: data = 8'hf5;
      17'd60712: data = 8'hf6;
      17'd60713: data = 8'hf5;
      17'd60714: data = 8'hf4;
      17'd60715: data = 8'hf4;
      17'd60716: data = 8'hf4;
      17'd60717: data = 8'hf5;
      17'd60718: data = 8'hf4;
      17'd60719: data = 8'hf5;
      17'd60720: data = 8'hf4;
      17'd60721: data = 8'hf5;
      17'd60722: data = 8'hf6;
      17'd60723: data = 8'hf9;
      17'd60724: data = 8'hf9;
      17'd60725: data = 8'hf5;
      17'd60726: data = 8'hf5;
      17'd60727: data = 8'hf5;
      17'd60728: data = 8'hf2;
      17'd60729: data = 8'hf2;
      17'd60730: data = 8'hf4;
      17'd60731: data = 8'hf4;
      17'd60732: data = 8'hf9;
      17'd60733: data = 8'hfa;
      17'd60734: data = 8'hfd;
      17'd60735: data = 8'hfe;
      17'd60736: data = 8'hfc;
      17'd60737: data = 8'hf6;
      17'd60738: data = 8'hf1;
      17'd60739: data = 8'hf2;
      17'd60740: data = 8'hf9;
      17'd60741: data = 8'hfa;
      17'd60742: data = 8'hf4;
      17'd60743: data = 8'hf2;
      17'd60744: data = 8'hf6;
      17'd60745: data = 8'hfc;
      17'd60746: data = 8'hfa;
      17'd60747: data = 8'hf2;
      17'd60748: data = 8'hf5;
      17'd60749: data = 8'hfa;
      17'd60750: data = 8'h01;
      17'd60751: data = 8'h05;
      17'd60752: data = 8'h00;
      17'd60753: data = 8'hfa;
      17'd60754: data = 8'h00;
      17'd60755: data = 8'h04;
      17'd60756: data = 8'h01;
      17'd60757: data = 8'h00;
      17'd60758: data = 8'h01;
      17'd60759: data = 8'h02;
      17'd60760: data = 8'h01;
      17'd60761: data = 8'h01;
      17'd60762: data = 8'hfc;
      17'd60763: data = 8'hf9;
      17'd60764: data = 8'hfc;
      17'd60765: data = 8'hfd;
      17'd60766: data = 8'hfd;
      17'd60767: data = 8'hfc;
      17'd60768: data = 8'hfc;
      17'd60769: data = 8'hfc;
      17'd60770: data = 8'hfc;
      17'd60771: data = 8'hfe;
      17'd60772: data = 8'h00;
      17'd60773: data = 8'hfc;
      17'd60774: data = 8'hf9;
      17'd60775: data = 8'hfa;
      17'd60776: data = 8'hfd;
      17'd60777: data = 8'h00;
      17'd60778: data = 8'hfc;
      17'd60779: data = 8'h00;
      17'd60780: data = 8'h05;
      17'd60781: data = 8'h06;
      17'd60782: data = 8'h01;
      17'd60783: data = 8'hfd;
      17'd60784: data = 8'h01;
      17'd60785: data = 8'h0a;
      17'd60786: data = 8'h02;
      17'd60787: data = 8'hfd;
      17'd60788: data = 8'h01;
      17'd60789: data = 8'hfc;
      17'd60790: data = 8'hf9;
      17'd60791: data = 8'hf9;
      17'd60792: data = 8'hf9;
      17'd60793: data = 8'hfc;
      17'd60794: data = 8'hf5;
      17'd60795: data = 8'hf9;
      17'd60796: data = 8'hfc;
      17'd60797: data = 8'hf4;
      17'd60798: data = 8'hf5;
      17'd60799: data = 8'hfe;
      17'd60800: data = 8'hfd;
      17'd60801: data = 8'hf9;
      17'd60802: data = 8'hf9;
      17'd60803: data = 8'h00;
      17'd60804: data = 8'h01;
      17'd60805: data = 8'hf9;
      17'd60806: data = 8'hfe;
      17'd60807: data = 8'h02;
      17'd60808: data = 8'h00;
      17'd60809: data = 8'hfe;
      17'd60810: data = 8'hfe;
      17'd60811: data = 8'hfe;
      17'd60812: data = 8'hfe;
      17'd60813: data = 8'hfc;
      17'd60814: data = 8'hfe;
      17'd60815: data = 8'h00;
      17'd60816: data = 8'hfd;
      17'd60817: data = 8'hfc;
      17'd60818: data = 8'hfd;
      17'd60819: data = 8'hfd;
      17'd60820: data = 8'hfc;
      17'd60821: data = 8'h00;
      17'd60822: data = 8'h00;
      17'd60823: data = 8'hfe;
      17'd60824: data = 8'hfe;
      17'd60825: data = 8'h01;
      17'd60826: data = 8'h04;
      17'd60827: data = 8'h01;
      17'd60828: data = 8'h02;
      17'd60829: data = 8'h05;
      17'd60830: data = 8'h0a;
      17'd60831: data = 8'h05;
      17'd60832: data = 8'h05;
      17'd60833: data = 8'h0a;
      17'd60834: data = 8'h09;
      17'd60835: data = 8'h0a;
      17'd60836: data = 8'h06;
      17'd60837: data = 8'h09;
      17'd60838: data = 8'h09;
      17'd60839: data = 8'h04;
      17'd60840: data = 8'h02;
      17'd60841: data = 8'h02;
      17'd60842: data = 8'h02;
      17'd60843: data = 8'h01;
      17'd60844: data = 8'h01;
      17'd60845: data = 8'h00;
      17'd60846: data = 8'h01;
      17'd60847: data = 8'h00;
      17'd60848: data = 8'h02;
      17'd60849: data = 8'h04;
      17'd60850: data = 8'h04;
      17'd60851: data = 8'h04;
      17'd60852: data = 8'h05;
      17'd60853: data = 8'h04;
      17'd60854: data = 8'h05;
      17'd60855: data = 8'h09;
      17'd60856: data = 8'h09;
      17'd60857: data = 8'h06;
      17'd60858: data = 8'h06;
      17'd60859: data = 8'h09;
      17'd60860: data = 8'h09;
      17'd60861: data = 8'h0a;
      17'd60862: data = 8'h09;
      17'd60863: data = 8'h0a;
      17'd60864: data = 8'h0d;
      17'd60865: data = 8'h0d;
      17'd60866: data = 8'h09;
      17'd60867: data = 8'h06;
      17'd60868: data = 8'h06;
      17'd60869: data = 8'h05;
      17'd60870: data = 8'h05;
      17'd60871: data = 8'h06;
      17'd60872: data = 8'h09;
      17'd60873: data = 8'h06;
      17'd60874: data = 8'h05;
      17'd60875: data = 8'h06;
      17'd60876: data = 8'h09;
      17'd60877: data = 8'h06;
      17'd60878: data = 8'h06;
      17'd60879: data = 8'h0a;
      17'd60880: data = 8'h0a;
      17'd60881: data = 8'h0a;
      17'd60882: data = 8'h09;
      17'd60883: data = 8'h09;
      17'd60884: data = 8'h09;
      17'd60885: data = 8'h09;
      17'd60886: data = 8'h09;
      17'd60887: data = 8'h09;
      17'd60888: data = 8'h05;
      17'd60889: data = 8'h02;
      17'd60890: data = 8'h04;
      17'd60891: data = 8'h02;
      17'd60892: data = 8'h02;
      17'd60893: data = 8'h01;
      17'd60894: data = 8'h02;
      17'd60895: data = 8'h02;
      17'd60896: data = 8'h02;
      17'd60897: data = 8'h01;
      17'd60898: data = 8'h01;
      17'd60899: data = 8'h00;
      17'd60900: data = 8'h01;
      17'd60901: data = 8'hfe;
      17'd60902: data = 8'hfc;
      17'd60903: data = 8'hfd;
      17'd60904: data = 8'hfa;
      17'd60905: data = 8'hfc;
      17'd60906: data = 8'h00;
      17'd60907: data = 8'h00;
      17'd60908: data = 8'h00;
      17'd60909: data = 8'h01;
      17'd60910: data = 8'h00;
      17'd60911: data = 8'h01;
      17'd60912: data = 8'h02;
      17'd60913: data = 8'hfe;
      17'd60914: data = 8'hfa;
      17'd60915: data = 8'hfc;
      17'd60916: data = 8'hfd;
      17'd60917: data = 8'h00;
      17'd60918: data = 8'h00;
      17'd60919: data = 8'hfa;
      17'd60920: data = 8'hf6;
      17'd60921: data = 8'hfa;
      17'd60922: data = 8'h00;
      17'd60923: data = 8'h01;
      17'd60924: data = 8'hfd;
      17'd60925: data = 8'hfa;
      17'd60926: data = 8'hfd;
      17'd60927: data = 8'h01;
      17'd60928: data = 8'h01;
      17'd60929: data = 8'hfe;
      17'd60930: data = 8'hfa;
      17'd60931: data = 8'hfd;
      17'd60932: data = 8'h00;
      17'd60933: data = 8'h00;
      17'd60934: data = 8'hfd;
      17'd60935: data = 8'hfc;
      17'd60936: data = 8'hfd;
      17'd60937: data = 8'h00;
      17'd60938: data = 8'h00;
      17'd60939: data = 8'hfd;
      17'd60940: data = 8'hf9;
      17'd60941: data = 8'hfc;
      17'd60942: data = 8'h00;
      17'd60943: data = 8'h01;
      17'd60944: data = 8'hfe;
      17'd60945: data = 8'hfd;
      17'd60946: data = 8'hfc;
      17'd60947: data = 8'hfc;
      17'd60948: data = 8'hfe;
      17'd60949: data = 8'hfa;
      17'd60950: data = 8'hfd;
      17'd60951: data = 8'hfe;
      17'd60952: data = 8'hfd;
      17'd60953: data = 8'hfd;
      17'd60954: data = 8'hfe;
      17'd60955: data = 8'hfe;
      17'd60956: data = 8'hfd;
      17'd60957: data = 8'hfd;
      17'd60958: data = 8'hfd;
      17'd60959: data = 8'hfe;
      17'd60960: data = 8'hfe;
      17'd60961: data = 8'hfd;
      17'd60962: data = 8'hfa;
      17'd60963: data = 8'hfe;
      17'd60964: data = 8'hfe;
      17'd60965: data = 8'h00;
      17'd60966: data = 8'h01;
      17'd60967: data = 8'h00;
      17'd60968: data = 8'h00;
      17'd60969: data = 8'hfe;
      17'd60970: data = 8'hfe;
      17'd60971: data = 8'hfd;
      17'd60972: data = 8'hfa;
      17'd60973: data = 8'hfa;
      17'd60974: data = 8'hfd;
      17'd60975: data = 8'hfd;
      17'd60976: data = 8'hfd;
      17'd60977: data = 8'hfa;
      17'd60978: data = 8'hfa;
      17'd60979: data = 8'hfd;
      17'd60980: data = 8'hfd;
      17'd60981: data = 8'hfc;
      17'd60982: data = 8'hfa;
      17'd60983: data = 8'hf9;
      17'd60984: data = 8'hfa;
      17'd60985: data = 8'hf9;
      17'd60986: data = 8'hf9;
      17'd60987: data = 8'hf6;
      17'd60988: data = 8'hf9;
      17'd60989: data = 8'hfe;
      17'd60990: data = 8'hfe;
      17'd60991: data = 8'h01;
      17'd60992: data = 8'hda;
      17'd60993: data = 8'hed;
      17'd60994: data = 8'h01;
      17'd60995: data = 8'he7;
      17'd60996: data = 8'hfa;
      17'd60997: data = 8'h06;
      17'd60998: data = 8'h01;
      17'd60999: data = 8'hf9;
      17'd61000: data = 8'h06;
      17'd61001: data = 8'h0a;
      17'd61002: data = 8'hfe;
      17'd61003: data = 8'hfd;
      17'd61004: data = 8'h01;
      17'd61005: data = 8'hec;
      17'd61006: data = 8'he7;
      17'd61007: data = 8'hf6;
      17'd61008: data = 8'hf1;
      17'd61009: data = 8'hec;
      17'd61010: data = 8'hf6;
      17'd61011: data = 8'hfd;
      17'd61012: data = 8'hf5;
      17'd61013: data = 8'hfc;
      17'd61014: data = 8'h06;
      17'd61015: data = 8'h04;
      17'd61016: data = 8'hfc;
      17'd61017: data = 8'h02;
      17'd61018: data = 8'h04;
      17'd61019: data = 8'hf6;
      17'd61020: data = 8'hfc;
      17'd61021: data = 8'hfc;
      17'd61022: data = 8'hec;
      17'd61023: data = 8'hf2;
      17'd61024: data = 8'hf6;
      17'd61025: data = 8'hf4;
      17'd61026: data = 8'hfc;
      17'd61027: data = 8'hf5;
      17'd61028: data = 8'h00;
      17'd61029: data = 8'h05;
      17'd61030: data = 8'h01;
      17'd61031: data = 8'h06;
      17'd61032: data = 8'h06;
      17'd61033: data = 8'h0c;
      17'd61034: data = 8'h0a;
      17'd61035: data = 8'hf4;
      17'd61036: data = 8'he9;
      17'd61037: data = 8'hf1;
      17'd61038: data = 8'heb;
      17'd61039: data = 8'hf2;
      17'd61040: data = 8'hfa;
      17'd61041: data = 8'h02;
      17'd61042: data = 8'h00;
      17'd61043: data = 8'h05;
      17'd61044: data = 8'h1a;
      17'd61045: data = 8'h1b;
      17'd61046: data = 8'h16;
      17'd61047: data = 8'h22;
      17'd61048: data = 8'h0e;
      17'd61049: data = 8'h04;
      17'd61050: data = 8'hfc;
      17'd61051: data = 8'he7;
      17'd61052: data = 8'he4;
      17'd61053: data = 8'hd1;
      17'd61054: data = 8'hde;
      17'd61055: data = 8'hf2;
      17'd61056: data = 8'hf4;
      17'd61057: data = 8'h0d;
      17'd61058: data = 8'h26;
      17'd61059: data = 8'h1f;
      17'd61060: data = 8'h24;
      17'd61061: data = 8'h27;
      17'd61062: data = 8'h24;
      17'd61063: data = 8'h12;
      17'd61064: data = 8'h04;
      17'd61065: data = 8'hef;
      17'd61066: data = 8'hda;
      17'd61067: data = 8'hd2;
      17'd61068: data = 8'hda;
      17'd61069: data = 8'he2;
      17'd61070: data = 8'he4;
      17'd61071: data = 8'hf5;
      17'd61072: data = 8'h05;
      17'd61073: data = 8'h0d;
      17'd61074: data = 8'h1a;
      17'd61075: data = 8'h24;
      17'd61076: data = 8'h23;
      17'd61077: data = 8'h22;
      17'd61078: data = 8'h0c;
      17'd61079: data = 8'h06;
      17'd61080: data = 8'hf1;
      17'd61081: data = 8'he5;
      17'd61082: data = 8'he2;
      17'd61083: data = 8'hde;
      17'd61084: data = 8'he9;
      17'd61085: data = 8'hf4;
      17'd61086: data = 8'hf6;
      17'd61087: data = 8'h00;
      17'd61088: data = 8'h05;
      17'd61089: data = 8'h16;
      17'd61090: data = 8'h15;
      17'd61091: data = 8'h0c;
      17'd61092: data = 8'h1a;
      17'd61093: data = 8'h0c;
      17'd61094: data = 8'h05;
      17'd61095: data = 8'h05;
      17'd61096: data = 8'h06;
      17'd61097: data = 8'hfa;
      17'd61098: data = 8'hfc;
      17'd61099: data = 8'h01;
      17'd61100: data = 8'h02;
      17'd61101: data = 8'h04;
      17'd61102: data = 8'h0c;
      17'd61103: data = 8'h0a;
      17'd61104: data = 8'h0c;
      17'd61105: data = 8'h0a;
      17'd61106: data = 8'h11;
      17'd61107: data = 8'h0d;
      17'd61108: data = 8'h05;
      17'd61109: data = 8'h09;
      17'd61110: data = 8'hfc;
      17'd61111: data = 8'hfa;
      17'd61112: data = 8'hf5;
      17'd61113: data = 8'hfa;
      17'd61114: data = 8'hf6;
      17'd61115: data = 8'hf4;
      17'd61116: data = 8'hf4;
      17'd61117: data = 8'h0a;
      17'd61118: data = 8'h00;
      17'd61119: data = 8'h12;
      17'd61120: data = 8'h11;
      17'd61121: data = 8'h06;
      17'd61122: data = 8'h0a;
      17'd61123: data = 8'h01;
      17'd61124: data = 8'h09;
      17'd61125: data = 8'hf5;
      17'd61126: data = 8'hf4;
      17'd61127: data = 8'hf5;
      17'd61128: data = 8'hf2;
      17'd61129: data = 8'hf6;
      17'd61130: data = 8'h02;
      17'd61131: data = 8'hf9;
      17'd61132: data = 8'h02;
      17'd61133: data = 8'h04;
      17'd61134: data = 8'h06;
      17'd61135: data = 8'h01;
      17'd61136: data = 8'h0c;
      17'd61137: data = 8'h06;
      17'd61138: data = 8'h06;
      17'd61139: data = 8'h0a;
      17'd61140: data = 8'hfd;
      17'd61141: data = 8'h0c;
      17'd61142: data = 8'hfc;
      17'd61143: data = 8'hf9;
      17'd61144: data = 8'h01;
      17'd61145: data = 8'hf6;
      17'd61146: data = 8'hf6;
      17'd61147: data = 8'h02;
      17'd61148: data = 8'h01;
      17'd61149: data = 8'h0d;
      17'd61150: data = 8'h05;
      17'd61151: data = 8'h00;
      17'd61152: data = 8'h06;
      17'd61153: data = 8'h04;
      17'd61154: data = 8'hf9;
      17'd61155: data = 8'h0c;
      17'd61156: data = 8'h01;
      17'd61157: data = 8'hfe;
      17'd61158: data = 8'hfa;
      17'd61159: data = 8'hef;
      17'd61160: data = 8'hfe;
      17'd61161: data = 8'hf9;
      17'd61162: data = 8'hfe;
      17'd61163: data = 8'hfc;
      17'd61164: data = 8'h02;
      17'd61165: data = 8'hf4;
      17'd61166: data = 8'hfd;
      17'd61167: data = 8'h02;
      17'd61168: data = 8'hfe;
      17'd61169: data = 8'h06;
      17'd61170: data = 8'h02;
      17'd61171: data = 8'h01;
      17'd61172: data = 8'h00;
      17'd61173: data = 8'hf5;
      17'd61174: data = 8'h00;
      17'd61175: data = 8'hef;
      17'd61176: data = 8'hed;
      17'd61177: data = 8'hfe;
      17'd61178: data = 8'hf4;
      17'd61179: data = 8'hfd;
      17'd61180: data = 8'hf9;
      17'd61181: data = 8'h01;
      17'd61182: data = 8'h01;
      17'd61183: data = 8'h04;
      17'd61184: data = 8'h02;
      17'd61185: data = 8'h09;
      17'd61186: data = 8'hfe;
      17'd61187: data = 8'hf9;
      17'd61188: data = 8'hfc;
      17'd61189: data = 8'hf5;
      17'd61190: data = 8'hf4;
      17'd61191: data = 8'h04;
      17'd61192: data = 8'hfe;
      17'd61193: data = 8'hf9;
      17'd61194: data = 8'h05;
      17'd61195: data = 8'hfc;
      17'd61196: data = 8'h05;
      17'd61197: data = 8'hf5;
      17'd61198: data = 8'h06;
      17'd61199: data = 8'h0a;
      17'd61200: data = 8'h0a;
      17'd61201: data = 8'h02;
      17'd61202: data = 8'hf6;
      17'd61203: data = 8'hfe;
      17'd61204: data = 8'hf6;
      17'd61205: data = 8'hf6;
      17'd61206: data = 8'heb;
      17'd61207: data = 8'hf6;
      17'd61208: data = 8'hed;
      17'd61209: data = 8'hf4;
      17'd61210: data = 8'h06;
      17'd61211: data = 8'h0a;
      17'd61212: data = 8'h15;
      17'd61213: data = 8'h19;
      17'd61214: data = 8'h13;
      17'd61215: data = 8'h22;
      17'd61216: data = 8'h12;
      17'd61217: data = 8'h15;
      17'd61218: data = 8'h04;
      17'd61219: data = 8'hfa;
      17'd61220: data = 8'hf1;
      17'd61221: data = 8'hf6;
      17'd61222: data = 8'hfa;
      17'd61223: data = 8'hed;
      17'd61224: data = 8'hfc;
      17'd61225: data = 8'hde;
      17'd61226: data = 8'h00;
      17'd61227: data = 8'hfe;
      17'd61228: data = 8'hfe;
      17'd61229: data = 8'h1c;
      17'd61230: data = 8'hfc;
      17'd61231: data = 8'hed;
      17'd61232: data = 8'hf1;
      17'd61233: data = 8'he7;
      17'd61234: data = 8'hf5;
      17'd61235: data = 8'he4;
      17'd61236: data = 8'he9;
      17'd61237: data = 8'he9;
      17'd61238: data = 8'he7;
      17'd61239: data = 8'h01;
      17'd61240: data = 8'h15;
      17'd61241: data = 8'h1c;
      17'd61242: data = 8'h1c;
      17'd61243: data = 8'h13;
      17'd61244: data = 8'h11;
      17'd61245: data = 8'h09;
      17'd61246: data = 8'hf9;
      17'd61247: data = 8'h00;
      17'd61248: data = 8'he7;
      17'd61249: data = 8'hd6;
      17'd61250: data = 8'he2;
      17'd61251: data = 8'hec;
      17'd61252: data = 8'heb;
      17'd61253: data = 8'h00;
      17'd61254: data = 8'hfd;
      17'd61255: data = 8'h04;
      17'd61256: data = 8'h06;
      17'd61257: data = 8'h0c;
      17'd61258: data = 8'h2c;
      17'd61259: data = 8'h12;
      17'd61260: data = 8'h11;
      17'd61261: data = 8'h26;
      17'd61262: data = 8'h04;
      17'd61263: data = 8'hf4;
      17'd61264: data = 8'hfa;
      17'd61265: data = 8'hec;
      17'd61266: data = 8'hec;
      17'd61267: data = 8'he5;
      17'd61268: data = 8'hf1;
      17'd61269: data = 8'h01;
      17'd61270: data = 8'hf1;
      17'd61271: data = 8'h02;
      17'd61272: data = 8'h1b;
      17'd61273: data = 8'h11;
      17'd61274: data = 8'h16;
      17'd61275: data = 8'h19;
      17'd61276: data = 8'h0a;
      17'd61277: data = 8'h0c;
      17'd61278: data = 8'hf9;
      17'd61279: data = 8'h01;
      17'd61280: data = 8'hfd;
      17'd61281: data = 8'he0;
      17'd61282: data = 8'hfc;
      17'd61283: data = 8'hf1;
      17'd61284: data = 8'he9;
      17'd61285: data = 8'hfc;
      17'd61286: data = 8'hfd;
      17'd61287: data = 8'h0a;
      17'd61288: data = 8'hfe;
      17'd61289: data = 8'h01;
      17'd61290: data = 8'h11;
      17'd61291: data = 8'h02;
      17'd61292: data = 8'hfe;
      17'd61293: data = 8'h04;
      17'd61294: data = 8'hfd;
      17'd61295: data = 8'he9;
      17'd61296: data = 8'heb;
      17'd61297: data = 8'hfe;
      17'd61298: data = 8'he7;
      17'd61299: data = 8'heb;
      17'd61300: data = 8'h0e;
      17'd61301: data = 8'h01;
      17'd61302: data = 8'h06;
      17'd61303: data = 8'h11;
      17'd61304: data = 8'h11;
      17'd61305: data = 8'h0a;
      17'd61306: data = 8'hfd;
      17'd61307: data = 8'h04;
      17'd61308: data = 8'hfc;
      17'd61309: data = 8'hfd;
      17'd61310: data = 8'hf4;
      17'd61311: data = 8'h00;
      17'd61312: data = 8'hfc;
      17'd61313: data = 8'hf9;
      17'd61314: data = 8'h09;
      17'd61315: data = 8'h0a;
      17'd61316: data = 8'h0e;
      17'd61317: data = 8'h12;
      17'd61318: data = 8'h1e;
      17'd61319: data = 8'h0a;
      17'd61320: data = 8'h0d;
      17'd61321: data = 8'h13;
      17'd61322: data = 8'h02;
      17'd61323: data = 8'h01;
      17'd61324: data = 8'hfd;
      17'd61325: data = 8'hfd;
      17'd61326: data = 8'hf1;
      17'd61327: data = 8'hec;
      17'd61328: data = 8'h00;
      17'd61329: data = 8'h00;
      17'd61330: data = 8'h01;
      17'd61331: data = 8'h01;
      17'd61332: data = 8'h0d;
      17'd61333: data = 8'h09;
      17'd61334: data = 8'h0c;
      17'd61335: data = 8'h0c;
      17'd61336: data = 8'h0a;
      17'd61337: data = 8'h05;
      17'd61338: data = 8'heb;
      17'd61339: data = 8'h02;
      17'd61340: data = 8'hfa;
      17'd61341: data = 8'hed;
      17'd61342: data = 8'hfc;
      17'd61343: data = 8'h00;
      17'd61344: data = 8'hed;
      17'd61345: data = 8'hf1;
      17'd61346: data = 8'h00;
      17'd61347: data = 8'h09;
      17'd61348: data = 8'hfd;
      17'd61349: data = 8'hf9;
      17'd61350: data = 8'h02;
      17'd61351: data = 8'hfd;
      17'd61352: data = 8'h00;
      17'd61353: data = 8'h05;
      17'd61354: data = 8'h15;
      17'd61355: data = 8'hfe;
      17'd61356: data = 8'h04;
      17'd61357: data = 8'h05;
      17'd61358: data = 8'hfd;
      17'd61359: data = 8'hfe;
      17'd61360: data = 8'hfa;
      17'd61361: data = 8'h05;
      17'd61362: data = 8'hf6;
      17'd61363: data = 8'hfc;
      17'd61364: data = 8'h04;
      17'd61365: data = 8'h04;
      17'd61366: data = 8'h01;
      17'd61367: data = 8'h02;
      17'd61368: data = 8'h00;
      17'd61369: data = 8'h00;
      17'd61370: data = 8'h04;
      17'd61371: data = 8'h02;
      17'd61372: data = 8'hf9;
      17'd61373: data = 8'hf9;
      17'd61374: data = 8'h00;
      17'd61375: data = 8'hf9;
      17'd61376: data = 8'hfe;
      17'd61377: data = 8'h04;
      17'd61378: data = 8'hfd;
      17'd61379: data = 8'hf2;
      17'd61380: data = 8'hf6;
      17'd61381: data = 8'h04;
      17'd61382: data = 8'hfe;
      17'd61383: data = 8'h01;
      17'd61384: data = 8'h02;
      17'd61385: data = 8'hf9;
      17'd61386: data = 8'hfc;
      17'd61387: data = 8'hfd;
      17'd61388: data = 8'h01;
      17'd61389: data = 8'hfd;
      17'd61390: data = 8'hf2;
      17'd61391: data = 8'hfc;
      17'd61392: data = 8'hf5;
      17'd61393: data = 8'hf2;
      17'd61394: data = 8'hfe;
      17'd61395: data = 8'hfd;
      17'd61396: data = 8'hef;
      17'd61397: data = 8'hf5;
      17'd61398: data = 8'hf5;
      17'd61399: data = 8'h01;
      17'd61400: data = 8'hfe;
      17'd61401: data = 8'hfa;
      17'd61402: data = 8'hfd;
      17'd61403: data = 8'hf1;
      17'd61404: data = 8'h01;
      17'd61405: data = 8'h09;
      17'd61406: data = 8'h05;
      17'd61407: data = 8'h04;
      17'd61408: data = 8'h02;
      17'd61409: data = 8'hf6;
      17'd61410: data = 8'h00;
      17'd61411: data = 8'h05;
      17'd61412: data = 8'h01;
      17'd61413: data = 8'h0c;
      17'd61414: data = 8'h05;
      17'd61415: data = 8'h13;
      17'd61416: data = 8'hef;
      17'd61417: data = 8'hd6;
      17'd61418: data = 8'hfe;
      17'd61419: data = 8'hf4;
      17'd61420: data = 8'he9;
      17'd61421: data = 8'hfd;
      17'd61422: data = 8'h01;
      17'd61423: data = 8'hfe;
      17'd61424: data = 8'hfe;
      17'd61425: data = 8'h11;
      17'd61426: data = 8'h12;
      17'd61427: data = 8'h00;
      17'd61428: data = 8'hf6;
      17'd61429: data = 8'h0a;
      17'd61430: data = 8'h02;
      17'd61431: data = 8'h01;
      17'd61432: data = 8'h0a;
      17'd61433: data = 8'h01;
      17'd61434: data = 8'h06;
      17'd61435: data = 8'hf4;
      17'd61436: data = 8'h0c;
      17'd61437: data = 8'h0c;
      17'd61438: data = 8'hfd;
      17'd61439: data = 8'h0a;
      17'd61440: data = 8'h09;
      17'd61441: data = 8'hfd;
      17'd61442: data = 8'hfd;
      17'd61443: data = 8'h0d;
      17'd61444: data = 8'h04;
      17'd61445: data = 8'hfa;
      17'd61446: data = 8'hed;
      17'd61447: data = 8'hf2;
      17'd61448: data = 8'hf4;
      17'd61449: data = 8'he7;
      17'd61450: data = 8'h04;
      17'd61451: data = 8'h0a;
      17'd61452: data = 8'hf2;
      17'd61453: data = 8'hfe;
      17'd61454: data = 8'h06;
      17'd61455: data = 8'h01;
      17'd61456: data = 8'hed;
      17'd61457: data = 8'hfd;
      17'd61458: data = 8'h02;
      17'd61459: data = 8'hf1;
      17'd61460: data = 8'hf1;
      17'd61461: data = 8'hf4;
      17'd61462: data = 8'hf9;
      17'd61463: data = 8'hef;
      17'd61464: data = 8'hf2;
      17'd61465: data = 8'hfe;
      17'd61466: data = 8'h05;
      17'd61467: data = 8'h06;
      17'd61468: data = 8'h01;
      17'd61469: data = 8'h05;
      17'd61470: data = 8'hf5;
      17'd61471: data = 8'hef;
      17'd61472: data = 8'hfd;
      17'd61473: data = 8'hfc;
      17'd61474: data = 8'h02;
      17'd61475: data = 8'h02;
      17'd61476: data = 8'hf9;
      17'd61477: data = 8'hfe;
      17'd61478: data = 8'h01;
      17'd61479: data = 8'h09;
      17'd61480: data = 8'h16;
      17'd61481: data = 8'h0d;
      17'd61482: data = 8'h0d;
      17'd61483: data = 8'h11;
      17'd61484: data = 8'h11;
      17'd61485: data = 8'h06;
      17'd61486: data = 8'h1a;
      17'd61487: data = 8'h15;
      17'd61488: data = 8'h00;
      17'd61489: data = 8'hfd;
      17'd61490: data = 8'hf9;
      17'd61491: data = 8'h04;
      17'd61492: data = 8'hfa;
      17'd61493: data = 8'hf4;
      17'd61494: data = 8'h06;
      17'd61495: data = 8'h02;
      17'd61496: data = 8'h05;
      17'd61497: data = 8'h05;
      17'd61498: data = 8'h0d;
      17'd61499: data = 8'hfc;
      17'd61500: data = 8'hec;
      17'd61501: data = 8'hfc;
      17'd61502: data = 8'he9;
      17'd61503: data = 8'he5;
      17'd61504: data = 8'he9;
      17'd61505: data = 8'hf1;
      17'd61506: data = 8'hed;
      17'd61507: data = 8'hfa;
      17'd61508: data = 8'h00;
      17'd61509: data = 8'h00;
      17'd61510: data = 8'h02;
      17'd61511: data = 8'hfc;
      17'd61512: data = 8'h05;
      17'd61513: data = 8'h09;
      17'd61514: data = 8'hfa;
      17'd61515: data = 8'h05;
      17'd61516: data = 8'h01;
      17'd61517: data = 8'hf2;
      17'd61518: data = 8'hf9;
      17'd61519: data = 8'hf6;
      17'd61520: data = 8'hf1;
      17'd61521: data = 8'hef;
      17'd61522: data = 8'hf9;
      17'd61523: data = 8'hfe;
      17'd61524: data = 8'hfc;
      17'd61525: data = 8'h06;
      17'd61526: data = 8'h12;
      17'd61527: data = 8'h0a;
      17'd61528: data = 8'h0c;
      17'd61529: data = 8'h11;
      17'd61530: data = 8'h0a;
      17'd61531: data = 8'h01;
      17'd61532: data = 8'hfa;
      17'd61533: data = 8'hf5;
      17'd61534: data = 8'hf2;
      17'd61535: data = 8'hf5;
      17'd61536: data = 8'hfd;
      17'd61537: data = 8'h02;
      17'd61538: data = 8'h01;
      17'd61539: data = 8'h05;
      17'd61540: data = 8'h09;
      17'd61541: data = 8'h06;
      17'd61542: data = 8'h0a;
      17'd61543: data = 8'h0a;
      17'd61544: data = 8'h06;
      17'd61545: data = 8'h00;
      17'd61546: data = 8'h06;
      17'd61547: data = 8'h06;
      17'd61548: data = 8'hfd;
      17'd61549: data = 8'h06;
      17'd61550: data = 8'h01;
      17'd61551: data = 8'hf1;
      17'd61552: data = 8'hfc;
      17'd61553: data = 8'h00;
      17'd61554: data = 8'hfc;
      17'd61555: data = 8'h04;
      17'd61556: data = 8'h09;
      17'd61557: data = 8'h04;
      17'd61558: data = 8'h0a;
      17'd61559: data = 8'h0e;
      17'd61560: data = 8'h12;
      17'd61561: data = 8'h0a;
      17'd61562: data = 8'h05;
      17'd61563: data = 8'h06;
      17'd61564: data = 8'h05;
      17'd61565: data = 8'h05;
      17'd61566: data = 8'h02;
      17'd61567: data = 8'h01;
      17'd61568: data = 8'h04;
      17'd61569: data = 8'hfd;
      17'd61570: data = 8'hf6;
      17'd61571: data = 8'hf4;
      17'd61572: data = 8'hf6;
      17'd61573: data = 8'hfa;
      17'd61574: data = 8'hf5;
      17'd61575: data = 8'hf5;
      17'd61576: data = 8'h02;
      17'd61577: data = 8'h09;
      17'd61578: data = 8'h0a;
      17'd61579: data = 8'h13;
      17'd61580: data = 8'h0c;
      17'd61581: data = 8'h05;
      17'd61582: data = 8'hfc;
      17'd61583: data = 8'hfc;
      17'd61584: data = 8'hfe;
      17'd61585: data = 8'hfd;
      17'd61586: data = 8'hf9;
      17'd61587: data = 8'hed;
      17'd61588: data = 8'hf1;
      17'd61589: data = 8'hf9;
      17'd61590: data = 8'hf9;
      17'd61591: data = 8'hfe;
      17'd61592: data = 8'h05;
      17'd61593: data = 8'h00;
      17'd61594: data = 8'h00;
      17'd61595: data = 8'h0c;
      17'd61596: data = 8'h0d;
      17'd61597: data = 8'h0a;
      17'd61598: data = 8'h0d;
      17'd61599: data = 8'h09;
      17'd61600: data = 8'h02;
      17'd61601: data = 8'hfd;
      17'd61602: data = 8'hfe;
      17'd61603: data = 8'h05;
      17'd61604: data = 8'hec;
      17'd61605: data = 8'hec;
      17'd61606: data = 8'h02;
      17'd61607: data = 8'hf6;
      17'd61608: data = 8'hfd;
      17'd61609: data = 8'h0d;
      17'd61610: data = 8'h0c;
      17'd61611: data = 8'h06;
      17'd61612: data = 8'h05;
      17'd61613: data = 8'h0e;
      17'd61614: data = 8'h0d;
      17'd61615: data = 8'h00;
      17'd61616: data = 8'hfe;
      17'd61617: data = 8'h00;
      17'd61618: data = 8'hf2;
      17'd61619: data = 8'hf1;
      17'd61620: data = 8'h00;
      17'd61621: data = 8'hfa;
      17'd61622: data = 8'hf1;
      17'd61623: data = 8'hf9;
      17'd61624: data = 8'hfc;
      17'd61625: data = 8'hf2;
      17'd61626: data = 8'hfa;
      17'd61627: data = 8'h05;
      17'd61628: data = 8'h04;
      17'd61629: data = 8'h00;
      17'd61630: data = 8'h01;
      17'd61631: data = 8'h04;
      17'd61632: data = 8'h02;
      17'd61633: data = 8'hf5;
      17'd61634: data = 8'hf5;
      17'd61635: data = 8'hf2;
      17'd61636: data = 8'he7;
      17'd61637: data = 8'hf6;
      17'd61638: data = 8'hf4;
      17'd61639: data = 8'hf2;
      17'd61640: data = 8'h00;
      17'd61641: data = 8'h01;
      17'd61642: data = 8'h02;
      17'd61643: data = 8'h05;
      17'd61644: data = 8'h04;
      17'd61645: data = 8'h0d;
      17'd61646: data = 8'h09;
      17'd61647: data = 8'hfc;
      17'd61648: data = 8'hfc;
      17'd61649: data = 8'hf9;
      17'd61650: data = 8'hf4;
      17'd61651: data = 8'hfc;
      17'd61652: data = 8'hfc;
      17'd61653: data = 8'hf9;
      17'd61654: data = 8'hf5;
      17'd61655: data = 8'hf6;
      17'd61656: data = 8'hfe;
      17'd61657: data = 8'h00;
      17'd61658: data = 8'h06;
      17'd61659: data = 8'h11;
      17'd61660: data = 8'h0a;
      17'd61661: data = 8'h04;
      17'd61662: data = 8'h0e;
      17'd61663: data = 8'h11;
      17'd61664: data = 8'h09;
      17'd61665: data = 8'hfe;
      17'd61666: data = 8'hfe;
      17'd61667: data = 8'hf6;
      17'd61668: data = 8'heb;
      17'd61669: data = 8'h00;
      17'd61670: data = 8'h05;
      17'd61671: data = 8'hf6;
      17'd61672: data = 8'hf4;
      17'd61673: data = 8'h02;
      17'd61674: data = 8'h04;
      17'd61675: data = 8'h04;
      17'd61676: data = 8'h12;
      17'd61677: data = 8'h11;
      17'd61678: data = 8'h00;
      17'd61679: data = 8'hf4;
      17'd61680: data = 8'h05;
      17'd61681: data = 8'h04;
      17'd61682: data = 8'hf4;
      17'd61683: data = 8'h00;
      17'd61684: data = 8'hf5;
      17'd61685: data = 8'hed;
      17'd61686: data = 8'hf6;
      17'd61687: data = 8'hfc;
      17'd61688: data = 8'hf9;
      17'd61689: data = 8'hf4;
      17'd61690: data = 8'hfd;
      17'd61691: data = 8'hfe;
      17'd61692: data = 8'h01;
      17'd61693: data = 8'h01;
      17'd61694: data = 8'h01;
      17'd61695: data = 8'hfc;
      17'd61696: data = 8'hf6;
      17'd61697: data = 8'hf9;
      17'd61698: data = 8'hf9;
      17'd61699: data = 8'hfe;
      17'd61700: data = 8'hf1;
      17'd61701: data = 8'hf2;
      17'd61702: data = 8'hfd;
      17'd61703: data = 8'hf6;
      17'd61704: data = 8'hfe;
      17'd61705: data = 8'h05;
      17'd61706: data = 8'hfa;
      17'd61707: data = 8'hfa;
      17'd61708: data = 8'hfd;
      17'd61709: data = 8'h00;
      17'd61710: data = 8'h04;
      17'd61711: data = 8'h05;
      17'd61712: data = 8'h04;
      17'd61713: data = 8'h04;
      17'd61714: data = 8'h05;
      17'd61715: data = 8'hfe;
      17'd61716: data = 8'h0c;
      17'd61717: data = 8'h01;
      17'd61718: data = 8'hfc;
      17'd61719: data = 8'h02;
      17'd61720: data = 8'hfe;
      17'd61721: data = 8'h01;
      17'd61722: data = 8'hfc;
      17'd61723: data = 8'h02;
      17'd61724: data = 8'h06;
      17'd61725: data = 8'hfd;
      17'd61726: data = 8'h00;
      17'd61727: data = 8'h01;
      17'd61728: data = 8'hfa;
      17'd61729: data = 8'h01;
      17'd61730: data = 8'h04;
      17'd61731: data = 8'h01;
      17'd61732: data = 8'h00;
      17'd61733: data = 8'hfc;
      17'd61734: data = 8'h05;
      17'd61735: data = 8'hfd;
      17'd61736: data = 8'hf2;
      17'd61737: data = 8'h02;
      17'd61738: data = 8'h02;
      17'd61739: data = 8'hf1;
      17'd61740: data = 8'hf1;
      17'd61741: data = 8'h00;
      17'd61742: data = 8'hef;
      17'd61743: data = 8'hf1;
      17'd61744: data = 8'hfd;
      17'd61745: data = 8'h04;
      17'd61746: data = 8'h04;
      17'd61747: data = 8'hfa;
      17'd61748: data = 8'h0a;
      17'd61749: data = 8'h00;
      17'd61750: data = 8'h05;
      17'd61751: data = 8'h0e;
      17'd61752: data = 8'hfe;
      17'd61753: data = 8'hfd;
      17'd61754: data = 8'hf9;
      17'd61755: data = 8'h05;
      17'd61756: data = 8'h02;
      17'd61757: data = 8'hf2;
      17'd61758: data = 8'hfe;
      17'd61759: data = 8'h05;
      17'd61760: data = 8'hfc;
      17'd61761: data = 8'h00;
      17'd61762: data = 8'h04;
      17'd61763: data = 8'h00;
      17'd61764: data = 8'h0e;
      17'd61765: data = 8'h0c;
      17'd61766: data = 8'h0c;
      17'd61767: data = 8'h0e;
      17'd61768: data = 8'h0c;
      17'd61769: data = 8'h06;
      17'd61770: data = 8'h00;
      17'd61771: data = 8'h01;
      17'd61772: data = 8'hfe;
      17'd61773: data = 8'h00;
      17'd61774: data = 8'h00;
      17'd61775: data = 8'h01;
      17'd61776: data = 8'h02;
      17'd61777: data = 8'h00;
      17'd61778: data = 8'h05;
      17'd61779: data = 8'h0e;
      17'd61780: data = 8'h0e;
      17'd61781: data = 8'h0d;
      17'd61782: data = 8'h05;
      17'd61783: data = 8'h05;
      17'd61784: data = 8'h06;
      17'd61785: data = 8'h00;
      17'd61786: data = 8'h01;
      17'd61787: data = 8'h01;
      17'd61788: data = 8'h00;
      17'd61789: data = 8'hf5;
      17'd61790: data = 8'hf4;
      17'd61791: data = 8'hfe;
      17'd61792: data = 8'hfe;
      17'd61793: data = 8'hfe;
      17'd61794: data = 8'h00;
      17'd61795: data = 8'h00;
      17'd61796: data = 8'h01;
      17'd61797: data = 8'h0a;
      17'd61798: data = 8'h11;
      17'd61799: data = 8'h02;
      17'd61800: data = 8'h02;
      17'd61801: data = 8'hf9;
      17'd61802: data = 8'hf4;
      17'd61803: data = 8'hf9;
      17'd61804: data = 8'hfe;
      17'd61805: data = 8'h00;
      17'd61806: data = 8'hec;
      17'd61807: data = 8'hf5;
      17'd61808: data = 8'h02;
      17'd61809: data = 8'h01;
      17'd61810: data = 8'h01;
      17'd61811: data = 8'h01;
      17'd61812: data = 8'h02;
      17'd61813: data = 8'hfe;
      17'd61814: data = 8'h00;
      17'd61815: data = 8'h02;
      17'd61816: data = 8'h02;
      17'd61817: data = 8'hfe;
      17'd61818: data = 8'hf9;
      17'd61819: data = 8'hfc;
      17'd61820: data = 8'hfa;
      17'd61821: data = 8'hfd;
      17'd61822: data = 8'h01;
      17'd61823: data = 8'h00;
      17'd61824: data = 8'hfe;
      17'd61825: data = 8'h00;
      17'd61826: data = 8'h02;
      17'd61827: data = 8'h00;
      17'd61828: data = 8'hfe;
      17'd61829: data = 8'h06;
      17'd61830: data = 8'h04;
      17'd61831: data = 8'hf6;
      17'd61832: data = 8'hf9;
      17'd61833: data = 8'hfd;
      17'd61834: data = 8'hfd;
      17'd61835: data = 8'hfe;
      17'd61836: data = 8'hfc;
      17'd61837: data = 8'hf5;
      17'd61838: data = 8'h02;
      17'd61839: data = 8'h0a;
      17'd61840: data = 8'h04;
      17'd61841: data = 8'h01;
      17'd61842: data = 8'hfd;
      17'd61843: data = 8'h00;
      17'd61844: data = 8'hfd;
      17'd61845: data = 8'hf6;
      17'd61846: data = 8'hf9;
      17'd61847: data = 8'hf5;
      17'd61848: data = 8'hf6;
      17'd61849: data = 8'hfa;
      17'd61850: data = 8'hfc;
      17'd61851: data = 8'hfc;
      17'd61852: data = 8'hf6;
      17'd61853: data = 8'hfa;
      17'd61854: data = 8'hfe;
      17'd61855: data = 8'h00;
      17'd61856: data = 8'h02;
      17'd61857: data = 8'h04;
      17'd61858: data = 8'h04;
      17'd61859: data = 8'h05;
      17'd61860: data = 8'h06;
      17'd61861: data = 8'h02;
      17'd61862: data = 8'hf9;
      17'd61863: data = 8'hf4;
      17'd61864: data = 8'hf5;
      17'd61865: data = 8'hf5;
      17'd61866: data = 8'hf4;
      17'd61867: data = 8'hf1;
      17'd61868: data = 8'hfc;
      17'd61869: data = 8'hfd;
      17'd61870: data = 8'hfc;
      17'd61871: data = 8'h04;
      17'd61872: data = 8'h00;
      17'd61873: data = 8'h02;
      17'd61874: data = 8'h04;
      17'd61875: data = 8'hfe;
      17'd61876: data = 8'hfd;
      17'd61877: data = 8'hfe;
      17'd61878: data = 8'h02;
      17'd61879: data = 8'h01;
      17'd61880: data = 8'hfd;
      17'd61881: data = 8'hfc;
      17'd61882: data = 8'hfc;
      17'd61883: data = 8'hfd;
      17'd61884: data = 8'hfd;
      17'd61885: data = 8'hfe;
      17'd61886: data = 8'hfc;
      17'd61887: data = 8'hfc;
      17'd61888: data = 8'hfe;
      17'd61889: data = 8'h00;
      17'd61890: data = 8'h09;
      17'd61891: data = 8'h04;
      17'd61892: data = 8'h04;
      17'd61893: data = 8'h04;
      17'd61894: data = 8'hfe;
      17'd61895: data = 8'h00;
      17'd61896: data = 8'h00;
      17'd61897: data = 8'h00;
      17'd61898: data = 8'hfd;
      17'd61899: data = 8'hfe;
      17'd61900: data = 8'h04;
      17'd61901: data = 8'h00;
      17'd61902: data = 8'hfe;
      17'd61903: data = 8'h01;
      17'd61904: data = 8'h01;
      17'd61905: data = 8'hfc;
      17'd61906: data = 8'hfc;
      17'd61907: data = 8'hfa;
      17'd61908: data = 8'hf6;
      17'd61909: data = 8'hf5;
      17'd61910: data = 8'hfc;
      17'd61911: data = 8'hfe;
      17'd61912: data = 8'hfa;
      17'd61913: data = 8'hfd;
      17'd61914: data = 8'hfc;
      17'd61915: data = 8'hfc;
      17'd61916: data = 8'hfc;
      17'd61917: data = 8'hfe;
      17'd61918: data = 8'h01;
      17'd61919: data = 8'hfd;
      17'd61920: data = 8'hfa;
      17'd61921: data = 8'h01;
      17'd61922: data = 8'h00;
      17'd61923: data = 8'hf9;
      17'd61924: data = 8'h00;
      17'd61925: data = 8'h01;
      17'd61926: data = 8'hfa;
      17'd61927: data = 8'hfc;
      17'd61928: data = 8'hfa;
      17'd61929: data = 8'h01;
      17'd61930: data = 8'h02;
      17'd61931: data = 8'h00;
      17'd61932: data = 8'h00;
      17'd61933: data = 8'h00;
      17'd61934: data = 8'h00;
      17'd61935: data = 8'h01;
      17'd61936: data = 8'h00;
      17'd61937: data = 8'hfd;
      17'd61938: data = 8'hf9;
      17'd61939: data = 8'hfc;
      17'd61940: data = 8'hfa;
      17'd61941: data = 8'hf5;
      17'd61942: data = 8'hfe;
      17'd61943: data = 8'h00;
      17'd61944: data = 8'hfe;
      17'd61945: data = 8'hfe;
      17'd61946: data = 8'h01;
      17'd61947: data = 8'h02;
      17'd61948: data = 8'h05;
      17'd61949: data = 8'h04;
      17'd61950: data = 8'hfd;
      17'd61951: data = 8'h01;
      17'd61952: data = 8'h0a;
      17'd61953: data = 8'h05;
      17'd61954: data = 8'h0a;
      17'd61955: data = 8'h04;
      17'd61956: data = 8'hfd;
      17'd61957: data = 8'h04;
      17'd61958: data = 8'h02;
      17'd61959: data = 8'h01;
      17'd61960: data = 8'h00;
      17'd61961: data = 8'hfc;
      17'd61962: data = 8'hfe;
      17'd61963: data = 8'h01;
      17'd61964: data = 8'h01;
      17'd61965: data = 8'h00;
      17'd61966: data = 8'hfe;
      17'd61967: data = 8'h00;
      17'd61968: data = 8'h04;
      17'd61969: data = 8'h01;
      17'd61970: data = 8'h04;
      17'd61971: data = 8'h09;
      17'd61972: data = 8'h01;
      17'd61973: data = 8'h00;
      17'd61974: data = 8'h05;
      17'd61975: data = 8'h04;
      17'd61976: data = 8'h02;
      17'd61977: data = 8'hfa;
      17'd61978: data = 8'hfd;
      17'd61979: data = 8'hfe;
      17'd61980: data = 8'hf4;
      17'd61981: data = 8'hfc;
      17'd61982: data = 8'hfa;
      17'd61983: data = 8'hfa;
      17'd61984: data = 8'h04;
      17'd61985: data = 8'hfe;
      17'd61986: data = 8'h04;
      17'd61987: data = 8'h02;
      17'd61988: data = 8'h05;
      17'd61989: data = 8'h15;
      17'd61990: data = 8'h06;
      17'd61991: data = 8'h01;
      17'd61992: data = 8'h04;
      17'd61993: data = 8'h01;
      17'd61994: data = 8'h01;
      17'd61995: data = 8'h00;
      17'd61996: data = 8'hfd;
      17'd61997: data = 8'hf9;
      17'd61998: data = 8'hf9;
      17'd61999: data = 8'hfd;
      17'd62000: data = 8'h00;
      17'd62001: data = 8'hfe;
      17'd62002: data = 8'hfe;
      17'd62003: data = 8'h02;
      17'd62004: data = 8'h06;
      17'd62005: data = 8'hfe;
      17'd62006: data = 8'h09;
      17'd62007: data = 8'h06;
      17'd62008: data = 8'h06;
      17'd62009: data = 8'h06;
      17'd62010: data = 8'hf9;
      17'd62011: data = 8'h00;
      17'd62012: data = 8'hfa;
      17'd62013: data = 8'hfe;
      17'd62014: data = 8'h02;
      17'd62015: data = 8'hfd;
      17'd62016: data = 8'h04;
      17'd62017: data = 8'h00;
      17'd62018: data = 8'h00;
      17'd62019: data = 8'h01;
      17'd62020: data = 8'h00;
      17'd62021: data = 8'h00;
      17'd62022: data = 8'hfe;
      17'd62023: data = 8'hfc;
      17'd62024: data = 8'hfe;
      17'd62025: data = 8'h00;
      17'd62026: data = 8'h02;
      17'd62027: data = 8'h04;
      17'd62028: data = 8'h00;
      17'd62029: data = 8'h00;
      17'd62030: data = 8'hfe;
      17'd62031: data = 8'hfe;
      17'd62032: data = 8'hfa;
      17'd62033: data = 8'hfa;
      17'd62034: data = 8'hfe;
      17'd62035: data = 8'hfc;
      17'd62036: data = 8'hfc;
      17'd62037: data = 8'hfe;
      17'd62038: data = 8'hfe;
      17'd62039: data = 8'hfa;
      17'd62040: data = 8'hfc;
      17'd62041: data = 8'hfc;
      17'd62042: data = 8'h00;
      17'd62043: data = 8'h09;
      17'd62044: data = 8'h05;
      17'd62045: data = 8'h01;
      17'd62046: data = 8'h02;
      17'd62047: data = 8'h04;
      17'd62048: data = 8'h05;
      17'd62049: data = 8'h00;
      17'd62050: data = 8'h02;
      17'd62051: data = 8'h02;
      17'd62052: data = 8'h00;
      17'd62053: data = 8'h00;
      17'd62054: data = 8'h01;
      17'd62055: data = 8'h04;
      17'd62056: data = 8'hfe;
      17'd62057: data = 8'hfe;
      17'd62058: data = 8'h00;
      17'd62059: data = 8'h00;
      17'd62060: data = 8'hfe;
      17'd62061: data = 8'h02;
      17'd62062: data = 8'h06;
      17'd62063: data = 8'h02;
      17'd62064: data = 8'h02;
      17'd62065: data = 8'h02;
      17'd62066: data = 8'h01;
      17'd62067: data = 8'h01;
      17'd62068: data = 8'h01;
      17'd62069: data = 8'hf6;
      17'd62070: data = 8'hed;
      17'd62071: data = 8'hed;
      17'd62072: data = 8'hf4;
      17'd62073: data = 8'hfd;
      17'd62074: data = 8'hfd;
      17'd62075: data = 8'h01;
      17'd62076: data = 8'h04;
      17'd62077: data = 8'h05;
      17'd62078: data = 8'h04;
      17'd62079: data = 8'h04;
      17'd62080: data = 8'h05;
      17'd62081: data = 8'h06;
      17'd62082: data = 8'h09;
      17'd62083: data = 8'h0a;
      17'd62084: data = 8'h05;
      17'd62085: data = 8'h06;
      17'd62086: data = 8'h11;
      17'd62087: data = 8'h0a;
      17'd62088: data = 8'h09;
      17'd62089: data = 8'h05;
      17'd62090: data = 8'hfe;
      17'd62091: data = 8'hf6;
      17'd62092: data = 8'hfc;
      17'd62093: data = 8'h00;
      17'd62094: data = 8'h00;
      17'd62095: data = 8'h01;
      17'd62096: data = 8'h04;
      17'd62097: data = 8'h06;
      17'd62098: data = 8'h09;
      17'd62099: data = 8'h05;
      17'd62100: data = 8'h01;
      17'd62101: data = 8'h01;
      17'd62102: data = 8'h01;
      17'd62103: data = 8'h02;
      17'd62104: data = 8'h00;
      17'd62105: data = 8'hfc;
      17'd62106: data = 8'hf9;
      17'd62107: data = 8'hfd;
      17'd62108: data = 8'hfa;
      17'd62109: data = 8'hfa;
      17'd62110: data = 8'hf5;
      17'd62111: data = 8'hf1;
      17'd62112: data = 8'hf1;
      17'd62113: data = 8'hef;
      17'd62114: data = 8'hed;
      17'd62115: data = 8'hed;
      17'd62116: data = 8'hf4;
      17'd62117: data = 8'hf4;
      17'd62118: data = 8'hef;
      17'd62119: data = 8'hf1;
      17'd62120: data = 8'hf1;
      17'd62121: data = 8'hf1;
      17'd62122: data = 8'hf1;
      17'd62123: data = 8'hf2;
      17'd62124: data = 8'hf5;
      17'd62125: data = 8'hf5;
      17'd62126: data = 8'hf5;
      17'd62127: data = 8'hf4;
      17'd62128: data = 8'hf6;
      17'd62129: data = 8'hf6;
      17'd62130: data = 8'hfa;
      17'd62131: data = 8'hfc;
      17'd62132: data = 8'hfe;
      17'd62133: data = 8'h01;
      17'd62134: data = 8'h00;
      17'd62135: data = 8'h01;
      17'd62136: data = 8'h05;
      17'd62137: data = 8'h05;
      17'd62138: data = 8'h06;
      17'd62139: data = 8'h0d;
      17'd62140: data = 8'h0d;
      17'd62141: data = 8'h0c;
      17'd62142: data = 8'h11;
      17'd62143: data = 8'h13;
      17'd62144: data = 8'h12;
      17'd62145: data = 8'h16;
      17'd62146: data = 8'h19;
      17'd62147: data = 8'h19;
      17'd62148: data = 8'h16;
      17'd62149: data = 8'h15;
      17'd62150: data = 8'h19;
      17'd62151: data = 8'h16;
      17'd62152: data = 8'h19;
      17'd62153: data = 8'h16;
      17'd62154: data = 8'h15;
      17'd62155: data = 8'h0e;
      17'd62156: data = 8'h0a;
      17'd62157: data = 8'h0a;
      17'd62158: data = 8'h05;
      17'd62159: data = 8'h04;
      17'd62160: data = 8'h02;
      17'd62161: data = 8'h01;
      17'd62162: data = 8'hfc;
      17'd62163: data = 8'hf9;
      17'd62164: data = 8'hf6;
      17'd62165: data = 8'hf4;
      17'd62166: data = 8'hf5;
      17'd62167: data = 8'hf4;
      17'd62168: data = 8'hf1;
      17'd62169: data = 8'hf2;
      17'd62170: data = 8'hf2;
      17'd62171: data = 8'hef;
      17'd62172: data = 8'hec;
      17'd62173: data = 8'hef;
      17'd62174: data = 8'hed;
      17'd62175: data = 8'hed;
      17'd62176: data = 8'hec;
      17'd62177: data = 8'heb;
      17'd62178: data = 8'hec;
      17'd62179: data = 8'hef;
      17'd62180: data = 8'hed;
      17'd62181: data = 8'hed;
      17'd62182: data = 8'hf1;
      17'd62183: data = 8'hef;
      17'd62184: data = 8'hf1;
      17'd62185: data = 8'hf4;
      17'd62186: data = 8'hf1;
      17'd62187: data = 8'hf2;
      17'd62188: data = 8'hf5;
      17'd62189: data = 8'hfa;
      17'd62190: data = 8'hf9;
      17'd62191: data = 8'hf9;
      17'd62192: data = 8'hfa;
      17'd62193: data = 8'hfa;
      17'd62194: data = 8'hfd;
      17'd62195: data = 8'hfe;
      17'd62196: data = 8'hfe;
      17'd62197: data = 8'hfd;
      17'd62198: data = 8'h00;
      17'd62199: data = 8'h01;
      17'd62200: data = 8'hfe;
      17'd62201: data = 8'h01;
      17'd62202: data = 8'h00;
      17'd62203: data = 8'hfd;
      17'd62204: data = 8'hfa;
      17'd62205: data = 8'hf9;
      17'd62206: data = 8'hfc;
      17'd62207: data = 8'hfd;
      17'd62208: data = 8'h00;
      17'd62209: data = 8'h00;
      17'd62210: data = 8'hfd;
      17'd62211: data = 8'hfa;
      17'd62212: data = 8'hfc;
      17'd62213: data = 8'hfe;
      17'd62214: data = 8'hfd;
      17'd62215: data = 8'hfa;
      17'd62216: data = 8'hf5;
      17'd62217: data = 8'hf6;
      17'd62218: data = 8'hf9;
      17'd62219: data = 8'hf9;
      17'd62220: data = 8'hf5;
      17'd62221: data = 8'hf2;
      17'd62222: data = 8'hf2;
      17'd62223: data = 8'hf4;
      17'd62224: data = 8'hf5;
      17'd62225: data = 8'hf4;
      17'd62226: data = 8'hf9;
      17'd62227: data = 8'hf4;
      17'd62228: data = 8'hf4;
      17'd62229: data = 8'hf4;
      17'd62230: data = 8'hf4;
      17'd62231: data = 8'hfa;
      17'd62232: data = 8'hf9;
      17'd62233: data = 8'hfc;
      17'd62234: data = 8'hfc;
      17'd62235: data = 8'hfa;
      17'd62236: data = 8'h00;
      17'd62237: data = 8'h02;
      17'd62238: data = 8'h02;
      17'd62239: data = 8'h02;
      17'd62240: data = 8'h09;
      17'd62241: data = 8'h06;
      17'd62242: data = 8'h0a;
      17'd62243: data = 8'h0c;
      17'd62244: data = 8'h0a;
      17'd62245: data = 8'h09;
      17'd62246: data = 8'h05;
      17'd62247: data = 8'h0c;
      17'd62248: data = 8'h0c;
      17'd62249: data = 8'h0c;
      17'd62250: data = 8'h0d;
      17'd62251: data = 8'h11;
      17'd62252: data = 8'h15;
      17'd62253: data = 8'h12;
      17'd62254: data = 8'h12;
      17'd62255: data = 8'h12;
      17'd62256: data = 8'h12;
      17'd62257: data = 8'h11;
      17'd62258: data = 8'h0d;
      17'd62259: data = 8'h0d;
      17'd62260: data = 8'h0e;
      17'd62261: data = 8'h0e;
      17'd62262: data = 8'h0c;
      17'd62263: data = 8'h0a;
      17'd62264: data = 8'h0a;
      17'd62265: data = 8'h0a;
      17'd62266: data = 8'h09;
      17'd62267: data = 8'h09;
      17'd62268: data = 8'h06;
      17'd62269: data = 8'h02;
      17'd62270: data = 8'h04;
      17'd62271: data = 8'h02;
      17'd62272: data = 8'h00;
      17'd62273: data = 8'h00;
      17'd62274: data = 8'h00;
      17'd62275: data = 8'h00;
      17'd62276: data = 8'h01;
      17'd62277: data = 8'h01;
      17'd62278: data = 8'h02;
      17'd62279: data = 8'h02;
      17'd62280: data = 8'h04;
      17'd62281: data = 8'h05;
      17'd62282: data = 8'h09;
      17'd62283: data = 8'h05;
      17'd62284: data = 8'h02;
      17'd62285: data = 8'h0a;
      17'd62286: data = 8'h06;
      17'd62287: data = 8'h05;
      17'd62288: data = 8'h05;
      17'd62289: data = 8'h02;
      17'd62290: data = 8'hfd;
      17'd62291: data = 8'hfc;
      17'd62292: data = 8'h00;
      17'd62293: data = 8'hfc;
      17'd62294: data = 8'h00;
      17'd62295: data = 8'h04;
      17'd62296: data = 8'h01;
      17'd62297: data = 8'h00;
      17'd62298: data = 8'h00;
      17'd62299: data = 8'hfc;
      17'd62300: data = 8'hfc;
      17'd62301: data = 8'hfa;
      17'd62302: data = 8'hfa;
      17'd62303: data = 8'h02;
      17'd62304: data = 8'h04;
      17'd62305: data = 8'h02;
      17'd62306: data = 8'h06;
      17'd62307: data = 8'h09;
      17'd62308: data = 8'h09;
      17'd62309: data = 8'h06;
      17'd62310: data = 8'h05;
      17'd62311: data = 8'h0a;
      17'd62312: data = 8'h0e;
      17'd62313: data = 8'h12;
      17'd62314: data = 8'h0a;
      17'd62315: data = 8'h12;
      17'd62316: data = 8'h16;
      17'd62317: data = 8'h13;
      17'd62318: data = 8'h12;
      17'd62319: data = 8'h0e;
      17'd62320: data = 8'h0a;
      17'd62321: data = 8'h06;
      17'd62322: data = 8'h06;
      17'd62323: data = 8'h06;
      17'd62324: data = 8'h06;
      17'd62325: data = 8'h05;
      17'd62326: data = 8'h09;
      17'd62327: data = 8'h05;
      17'd62328: data = 8'h00;
      17'd62329: data = 8'hfc;
      17'd62330: data = 8'h00;
      17'd62331: data = 8'h04;
      17'd62332: data = 8'hfc;
      17'd62333: data = 8'hfa;
      17'd62334: data = 8'h00;
      17'd62335: data = 8'hfe;
      17'd62336: data = 8'hfc;
      17'd62337: data = 8'hfc;
      17'd62338: data = 8'hfe;
      17'd62339: data = 8'hfe;
      17'd62340: data = 8'hfa;
      17'd62341: data = 8'hf5;
      17'd62342: data = 8'hef;
      17'd62343: data = 8'hec;
      17'd62344: data = 8'heb;
      17'd62345: data = 8'hed;
      17'd62346: data = 8'hed;
      17'd62347: data = 8'he9;
      17'd62348: data = 8'heb;
      17'd62349: data = 8'heb;
      17'd62350: data = 8'he7;
      17'd62351: data = 8'he5;
      17'd62352: data = 8'he9;
      17'd62353: data = 8'hec;
      17'd62354: data = 8'hec;
      17'd62355: data = 8'he7;
      17'd62356: data = 8'heb;
      17'd62357: data = 8'hed;
      17'd62358: data = 8'hf1;
      17'd62359: data = 8'hef;
      17'd62360: data = 8'hf2;
      17'd62361: data = 8'hf5;
      17'd62362: data = 8'hf5;
      17'd62363: data = 8'hfa;
      17'd62364: data = 8'hf9;
      17'd62365: data = 8'hfc;
      17'd62366: data = 8'h02;
      17'd62367: data = 8'h04;
      17'd62368: data = 8'h05;
      17'd62369: data = 8'h04;
      17'd62370: data = 8'h05;
      17'd62371: data = 8'h09;
      17'd62372: data = 8'h0a;
      17'd62373: data = 8'h06;
      17'd62374: data = 8'h04;
      17'd62375: data = 8'h09;
      17'd62376: data = 8'h0c;
      17'd62377: data = 8'h09;
      17'd62378: data = 8'h06;
      17'd62379: data = 8'h06;
      17'd62380: data = 8'h0c;
      17'd62381: data = 8'h0e;
      17'd62382: data = 8'h0d;
      17'd62383: data = 8'h0d;
      17'd62384: data = 8'h0d;
      17'd62385: data = 8'h0a;
      17'd62386: data = 8'h09;
      17'd62387: data = 8'h05;
      17'd62388: data = 8'h04;
      17'd62389: data = 8'h09;
      17'd62390: data = 8'h09;
      17'd62391: data = 8'h04;
      17'd62392: data = 8'hfe;
      17'd62393: data = 8'hfd;
      17'd62394: data = 8'hfe;
      17'd62395: data = 8'h00;
      17'd62396: data = 8'hfa;
      17'd62397: data = 8'hf5;
      17'd62398: data = 8'hf6;
      17'd62399: data = 8'hf6;
      17'd62400: data = 8'hf4;
      17'd62401: data = 8'hf1;
      17'd62402: data = 8'hef;
      17'd62403: data = 8'hf1;
      17'd62404: data = 8'hef;
      17'd62405: data = 8'hec;
      17'd62406: data = 8'heb;
      17'd62407: data = 8'heb;
      17'd62408: data = 8'heb;
      17'd62409: data = 8'hed;
      17'd62410: data = 8'hef;
      17'd62411: data = 8'hef;
      17'd62412: data = 8'hf1;
      17'd62413: data = 8'hf1;
      17'd62414: data = 8'hf1;
      17'd62415: data = 8'hed;
      17'd62416: data = 8'hed;
      17'd62417: data = 8'hf4;
      17'd62418: data = 8'hf4;
      17'd62419: data = 8'hf1;
      17'd62420: data = 8'hed;
      17'd62421: data = 8'hf2;
      17'd62422: data = 8'hf4;
      17'd62423: data = 8'hf5;
      17'd62424: data = 8'hf2;
      17'd62425: data = 8'hf2;
      17'd62426: data = 8'hf5;
      17'd62427: data = 8'hf4;
      17'd62428: data = 8'hf5;
      17'd62429: data = 8'hf5;
      17'd62430: data = 8'hf5;
      17'd62431: data = 8'hf5;
      17'd62432: data = 8'hf6;
      17'd62433: data = 8'hf6;
      17'd62434: data = 8'hf5;
      17'd62435: data = 8'hf5;
      17'd62436: data = 8'hf5;
      17'd62437: data = 8'hf5;
      17'd62438: data = 8'hf5;
      17'd62439: data = 8'hf4;
      17'd62440: data = 8'hf6;
      17'd62441: data = 8'hf9;
      17'd62442: data = 8'hf5;
      17'd62443: data = 8'hf5;
      17'd62444: data = 8'hf6;
      17'd62445: data = 8'hf6;
      17'd62446: data = 8'hf6;
      17'd62447: data = 8'hf9;
      17'd62448: data = 8'hf5;
      17'd62449: data = 8'hf9;
      17'd62450: data = 8'hfa;
      17'd62451: data = 8'hf9;
      17'd62452: data = 8'hf9;
      17'd62453: data = 8'hf9;
      17'd62454: data = 8'hf6;
      17'd62455: data = 8'hfa;
      17'd62456: data = 8'hf6;
      17'd62457: data = 8'hf5;
      17'd62458: data = 8'hf9;
      17'd62459: data = 8'hfa;
      17'd62460: data = 8'hfd;
      17'd62461: data = 8'hfe;
      17'd62462: data = 8'h00;
      17'd62463: data = 8'h01;
      17'd62464: data = 8'h02;
      17'd62465: data = 8'h00;
      17'd62466: data = 8'h02;
      17'd62467: data = 8'h02;
      17'd62468: data = 8'h02;
      17'd62469: data = 8'h04;
      17'd62470: data = 8'h01;
      17'd62471: data = 8'h05;
      17'd62472: data = 8'h05;
      17'd62473: data = 8'h06;
      17'd62474: data = 8'h06;
      17'd62475: data = 8'h09;
      17'd62476: data = 8'h0a;
      17'd62477: data = 8'h0d;
      17'd62478: data = 8'h0e;
      17'd62479: data = 8'h11;
      17'd62480: data = 8'h12;
      17'd62481: data = 8'h12;
      17'd62482: data = 8'h13;
      17'd62483: data = 8'h13;
      17'd62484: data = 8'h12;
      17'd62485: data = 8'h12;
      17'd62486: data = 8'h12;
      17'd62487: data = 8'h0e;
      17'd62488: data = 8'h11;
      17'd62489: data = 8'h12;
      17'd62490: data = 8'h13;
      17'd62491: data = 8'h13;
      17'd62492: data = 8'h13;
      17'd62493: data = 8'h12;
      17'd62494: data = 8'h12;
      17'd62495: data = 8'h12;
      17'd62496: data = 8'h13;
      17'd62497: data = 8'h16;
      17'd62498: data = 8'h13;
      17'd62499: data = 8'h12;
      17'd62500: data = 8'h11;
      17'd62501: data = 8'h11;
      17'd62502: data = 8'h11;
      17'd62503: data = 8'h12;
      17'd62504: data = 8'h11;
      17'd62505: data = 8'h12;
      17'd62506: data = 8'h15;
      17'd62507: data = 8'h11;
      17'd62508: data = 8'h11;
      17'd62509: data = 8'h12;
      17'd62510: data = 8'h16;
      17'd62511: data = 8'h15;
      17'd62512: data = 8'h11;
      17'd62513: data = 8'h0c;
      17'd62514: data = 8'h0c;
      17'd62515: data = 8'h0a;
      17'd62516: data = 8'h0a;
      17'd62517: data = 8'h0a;
      17'd62518: data = 8'h09;
      17'd62519: data = 8'h09;
      17'd62520: data = 8'h09;
      17'd62521: data = 8'h0a;
      17'd62522: data = 8'h0a;
      17'd62523: data = 8'h0a;
      17'd62524: data = 8'h06;
      17'd62525: data = 8'h06;
      17'd62526: data = 8'h09;
      17'd62527: data = 8'h04;
      17'd62528: data = 8'h05;
      17'd62529: data = 8'h05;
      17'd62530: data = 8'h02;
      17'd62531: data = 8'h01;
      17'd62532: data = 8'h01;
      17'd62533: data = 8'h01;
      17'd62534: data = 8'h00;
      17'd62535: data = 8'hfd;
      17'd62536: data = 8'hfc;
      17'd62537: data = 8'hfe;
      17'd62538: data = 8'h01;
      17'd62539: data = 8'hfe;
      17'd62540: data = 8'hfd;
      17'd62541: data = 8'hfe;
      17'd62542: data = 8'hfe;
      17'd62543: data = 8'h01;
      17'd62544: data = 8'h00;
      17'd62545: data = 8'hfa;
      17'd62546: data = 8'hf6;
      17'd62547: data = 8'hf6;
      17'd62548: data = 8'hfa;
      17'd62549: data = 8'hfd;
      17'd62550: data = 8'hfe;
      17'd62551: data = 8'hfd;
      17'd62552: data = 8'h00;
      17'd62553: data = 8'h06;
      17'd62554: data = 8'h09;
      17'd62555: data = 8'h00;
      17'd62556: data = 8'hfe;
      17'd62557: data = 8'h00;
      17'd62558: data = 8'h00;
      17'd62559: data = 8'hfe;
      17'd62560: data = 8'h01;
      17'd62561: data = 8'h01;
      17'd62562: data = 8'h01;
      17'd62563: data = 8'h04;
      17'd62564: data = 8'h02;
      17'd62565: data = 8'h04;
      17'd62566: data = 8'h00;
      17'd62567: data = 8'hfd;
      17'd62568: data = 8'hfe;
      17'd62569: data = 8'h02;
      17'd62570: data = 8'h01;
      17'd62571: data = 8'h01;
      17'd62572: data = 8'h05;
      17'd62573: data = 8'h02;
      17'd62574: data = 8'h01;
      17'd62575: data = 8'h02;
      17'd62576: data = 8'h01;
      17'd62577: data = 8'h00;
      17'd62578: data = 8'hfe;
      17'd62579: data = 8'hfc;
      17'd62580: data = 8'h00;
      17'd62581: data = 8'h02;
      17'd62582: data = 8'h00;
      17'd62583: data = 8'h02;
      17'd62584: data = 8'h05;
      17'd62585: data = 8'h04;
      17'd62586: data = 8'h02;
      17'd62587: data = 8'hfe;
      17'd62588: data = 8'hf9;
      17'd62589: data = 8'hf5;
      17'd62590: data = 8'hf5;
      17'd62591: data = 8'hf4;
      17'd62592: data = 8'hf2;
      17'd62593: data = 8'hf1;
      17'd62594: data = 8'hf2;
      17'd62595: data = 8'hf2;
      17'd62596: data = 8'hef;
      17'd62597: data = 8'hef;
      17'd62598: data = 8'hec;
      17'd62599: data = 8'hec;
      17'd62600: data = 8'hed;
      17'd62601: data = 8'hec;
      17'd62602: data = 8'hed;
      17'd62603: data = 8'hed;
      17'd62604: data = 8'hef;
      17'd62605: data = 8'hf1;
      17'd62606: data = 8'hed;
      17'd62607: data = 8'hed;
      17'd62608: data = 8'hec;
      17'd62609: data = 8'he7;
      17'd62610: data = 8'he4;
      17'd62611: data = 8'he7;
      17'd62612: data = 8'hec;
      17'd62613: data = 8'hed;
      17'd62614: data = 8'hef;
      17'd62615: data = 8'hf1;
      17'd62616: data = 8'hf4;
      17'd62617: data = 8'hf5;
      17'd62618: data = 8'hf2;
      17'd62619: data = 8'hec;
      17'd62620: data = 8'hec;
      17'd62621: data = 8'hec;
      17'd62622: data = 8'hec;
      17'd62623: data = 8'hef;
      17'd62624: data = 8'hf1;
      17'd62625: data = 8'hf5;
      17'd62626: data = 8'hf9;
      17'd62627: data = 8'hf9;
      17'd62628: data = 8'hfa;
      17'd62629: data = 8'hfd;
      17'd62630: data = 8'hfc;
      17'd62631: data = 8'hfd;
      17'd62632: data = 8'hfe;
      17'd62633: data = 8'hfe;
      17'd62634: data = 8'h00;
      17'd62635: data = 8'h01;
      17'd62636: data = 8'h01;
      17'd62637: data = 8'h01;
      17'd62638: data = 8'h01;
      17'd62639: data = 8'hfe;
      17'd62640: data = 8'hfd;
      17'd62641: data = 8'hfd;
      17'd62642: data = 8'hfe;
      17'd62643: data = 8'hfd;
      17'd62644: data = 8'h00;
      17'd62645: data = 8'h02;
      17'd62646: data = 8'h04;
      17'd62647: data = 8'h02;
      17'd62648: data = 8'h01;
      17'd62649: data = 8'h00;
      17'd62650: data = 8'h00;
      17'd62651: data = 8'hfe;
      17'd62652: data = 8'hfc;
      17'd62653: data = 8'hfd;
      17'd62654: data = 8'hfe;
      17'd62655: data = 8'hfd;
      17'd62656: data = 8'h00;
      17'd62657: data = 8'h00;
      17'd62658: data = 8'h01;
      17'd62659: data = 8'h02;
      17'd62660: data = 8'h01;
      17'd62661: data = 8'h02;
      17'd62662: data = 8'hfe;
      17'd62663: data = 8'h00;
      17'd62664: data = 8'h01;
      17'd62665: data = 8'h01;
      17'd62666: data = 8'hfd;
      17'd62667: data = 8'hfc;
      17'd62668: data = 8'h00;
      17'd62669: data = 8'hfa;
      17'd62670: data = 8'hf6;
      17'd62671: data = 8'hf6;
      17'd62672: data = 8'hfa;
      17'd62673: data = 8'hfc;
      17'd62674: data = 8'hfc;
      17'd62675: data = 8'hfd;
      17'd62676: data = 8'hfd;
      17'd62677: data = 8'h00;
      17'd62678: data = 8'h00;
      17'd62679: data = 8'hfd;
      17'd62680: data = 8'hfa;
      17'd62681: data = 8'hf6;
      17'd62682: data = 8'hfa;
      17'd62683: data = 8'hf6;
      17'd62684: data = 8'hf6;
      17'd62685: data = 8'hf9;
      17'd62686: data = 8'hf9;
      17'd62687: data = 8'hf5;
      17'd62688: data = 8'hf6;
      17'd62689: data = 8'hf9;
      17'd62690: data = 8'hf6;
      17'd62691: data = 8'hf5;
      17'd62692: data = 8'hf5;
      17'd62693: data = 8'hf2;
      17'd62694: data = 8'hf1;
      17'd62695: data = 8'hf1;
      17'd62696: data = 8'hf2;
      17'd62697: data = 8'hf5;
      17'd62698: data = 8'hf2;
      17'd62699: data = 8'hf1;
      17'd62700: data = 8'hf4;
      17'd62701: data = 8'hf5;
      17'd62702: data = 8'hf1;
      17'd62703: data = 8'hf2;
      17'd62704: data = 8'hf5;
      17'd62705: data = 8'hf5;
      17'd62706: data = 8'hf5;
      17'd62707: data = 8'hf5;
      17'd62708: data = 8'hf6;
      17'd62709: data = 8'hf9;
      17'd62710: data = 8'hf9;
      17'd62711: data = 8'hfa;
      17'd62712: data = 8'hfc;
      17'd62713: data = 8'hf5;
      17'd62714: data = 8'hf6;
      17'd62715: data = 8'hfc;
      17'd62716: data = 8'hfa;
      17'd62717: data = 8'hf9;
      17'd62718: data = 8'hfc;
      17'd62719: data = 8'hfe;
      17'd62720: data = 8'hfe;
      17'd62721: data = 8'h00;
      17'd62722: data = 8'hfe;
      17'd62723: data = 8'h01;
      17'd62724: data = 8'h04;
      17'd62725: data = 8'h04;
      17'd62726: data = 8'h02;
      17'd62727: data = 8'h01;
      17'd62728: data = 8'h04;
      17'd62729: data = 8'h0a;
      17'd62730: data = 8'h0c;
      17'd62731: data = 8'h0c;
      17'd62732: data = 8'h0d;
      17'd62733: data = 8'h0c;
      17'd62734: data = 8'h11;
      17'd62735: data = 8'h11;
      17'd62736: data = 8'h0e;
      17'd62737: data = 8'h0e;
      17'd62738: data = 8'h12;
      17'd62739: data = 8'h15;
      17'd62740: data = 8'h12;
      17'd62741: data = 8'h0d;
      17'd62742: data = 8'h0e;
      17'd62743: data = 8'h13;
      17'd62744: data = 8'h15;
      17'd62745: data = 8'h15;
      17'd62746: data = 8'h12;
      17'd62747: data = 8'h13;
      17'd62748: data = 8'h19;
      17'd62749: data = 8'h19;
      17'd62750: data = 8'h16;
      17'd62751: data = 8'h11;
      17'd62752: data = 8'h11;
      17'd62753: data = 8'h16;
      17'd62754: data = 8'h19;
      17'd62755: data = 8'h15;
      17'd62756: data = 8'h19;
      17'd62757: data = 8'h1a;
      17'd62758: data = 8'h19;
      17'd62759: data = 8'h16;
      17'd62760: data = 8'h12;
      17'd62761: data = 8'h15;
      17'd62762: data = 8'h1a;
      17'd62763: data = 8'h19;
      17'd62764: data = 8'h19;
      17'd62765: data = 8'h15;
      17'd62766: data = 8'h12;
      17'd62767: data = 8'h15;
      17'd62768: data = 8'h13;
      17'd62769: data = 8'h13;
      17'd62770: data = 8'h0e;
      17'd62771: data = 8'h0c;
      17'd62772: data = 8'h0c;
      17'd62773: data = 8'h0d;
      17'd62774: data = 8'h0e;
      17'd62775: data = 8'h0e;
      17'd62776: data = 8'h0e;
      17'd62777: data = 8'h0c;
      17'd62778: data = 8'h0a;
      17'd62779: data = 8'h0a;
      17'd62780: data = 8'h0a;
      17'd62781: data = 8'h0a;
      17'd62782: data = 8'h06;
      17'd62783: data = 8'h06;
      17'd62784: data = 8'h06;
      17'd62785: data = 8'h02;
      17'd62786: data = 8'h02;
      17'd62787: data = 8'h02;
      17'd62788: data = 8'hfe;
      17'd62789: data = 8'hfc;
      17'd62790: data = 8'hfe;
      17'd62791: data = 8'h00;
      17'd62792: data = 8'hfe;
      17'd62793: data = 8'hfd;
      17'd62794: data = 8'h00;
      17'd62795: data = 8'h01;
      17'd62796: data = 8'hfe;
      17'd62797: data = 8'hfa;
      17'd62798: data = 8'hfa;
      17'd62799: data = 8'hfe;
      17'd62800: data = 8'hfe;
      17'd62801: data = 8'hfa;
      17'd62802: data = 8'hf9;
      17'd62803: data = 8'hfa;
      17'd62804: data = 8'hfe;
      17'd62805: data = 8'hfe;
      17'd62806: data = 8'h00;
      17'd62807: data = 8'h01;
      17'd62808: data = 8'h01;
      17'd62809: data = 8'h01;
      17'd62810: data = 8'h00;
      17'd62811: data = 8'h00;
      17'd62812: data = 8'hfd;
      17'd62813: data = 8'h02;
      17'd62814: data = 8'h04;
      17'd62815: data = 8'h02;
      17'd62816: data = 8'h04;
      17'd62817: data = 8'h04;
      17'd62818: data = 8'h02;
      17'd62819: data = 8'h02;
      17'd62820: data = 8'h00;
      17'd62821: data = 8'hfe;
      17'd62822: data = 8'h02;
      17'd62823: data = 8'h05;
      17'd62824: data = 8'h04;
      17'd62825: data = 8'h04;
      17'd62826: data = 8'h06;
      17'd62827: data = 8'h06;
      17'd62828: data = 8'h05;
      17'd62829: data = 8'h01;
      17'd62830: data = 8'h00;
      17'd62831: data = 8'h00;
      17'd62832: data = 8'h00;
      17'd62833: data = 8'h00;
      17'd62834: data = 8'h00;
      17'd62835: data = 8'h02;
      17'd62836: data = 8'h04;
      17'd62837: data = 8'h02;
      17'd62838: data = 8'h01;
      17'd62839: data = 8'h00;
      17'd62840: data = 8'hfe;
      17'd62841: data = 8'hf9;
      17'd62842: data = 8'hf5;
      17'd62843: data = 8'hf9;
      17'd62844: data = 8'hf4;
      17'd62845: data = 8'hf2;
      17'd62846: data = 8'hf4;
      17'd62847: data = 8'hf4;
      17'd62848: data = 8'hf2;
      17'd62849: data = 8'hef;
      17'd62850: data = 8'hed;
      17'd62851: data = 8'hec;
      17'd62852: data = 8'hec;
      17'd62853: data = 8'hec;
      17'd62854: data = 8'hec;
      17'd62855: data = 8'hec;
      17'd62856: data = 8'heb;
      17'd62857: data = 8'heb;
      17'd62858: data = 8'heb;
      17'd62859: data = 8'he9;
      17'd62860: data = 8'he9;
      17'd62861: data = 8'he7;
      17'd62862: data = 8'he9;
      17'd62863: data = 8'he7;
      17'd62864: data = 8'he9;
      17'd62865: data = 8'heb;
      17'd62866: data = 8'hef;
      17'd62867: data = 8'hf1;
      17'd62868: data = 8'hef;
      17'd62869: data = 8'hf4;
      17'd62870: data = 8'hf2;
      17'd62871: data = 8'hf1;
      17'd62872: data = 8'hed;
      17'd62873: data = 8'hec;
      17'd62874: data = 8'hef;
      17'd62875: data = 8'hef;
      17'd62876: data = 8'hf1;
      17'd62877: data = 8'hf4;
      17'd62878: data = 8'hf5;
      17'd62879: data = 8'hfa;
      17'd62880: data = 8'hfa;
      17'd62881: data = 8'hfd;
      17'd62882: data = 8'hfc;
      17'd62883: data = 8'hfc;
      17'd62884: data = 8'hfa;
      17'd62885: data = 8'hf6;
      17'd62886: data = 8'hfa;
      17'd62887: data = 8'hfc;
      17'd62888: data = 8'hfe;
      17'd62889: data = 8'h00;
      17'd62890: data = 8'h00;
      17'd62891: data = 8'hfe;
      17'd62892: data = 8'hfd;
      17'd62893: data = 8'hfc;
      17'd62894: data = 8'hf6;
      17'd62895: data = 8'hfc;
      17'd62896: data = 8'hfd;
      17'd62897: data = 8'hfd;
      17'd62898: data = 8'h00;
      17'd62899: data = 8'h00;
      17'd62900: data = 8'h01;
      17'd62901: data = 8'h02;
      17'd62902: data = 8'h00;
      17'd62903: data = 8'h00;
      17'd62904: data = 8'h00;
      17'd62905: data = 8'h00;
      17'd62906: data = 8'hfe;
      17'd62907: data = 8'h00;
      17'd62908: data = 8'h02;
      17'd62909: data = 8'h04;
      17'd62910: data = 8'h04;
      17'd62911: data = 8'h02;
      17'd62912: data = 8'h02;
      17'd62913: data = 8'h02;
      17'd62914: data = 8'h02;
      17'd62915: data = 8'h04;
      17'd62916: data = 8'h04;
      17'd62917: data = 8'h00;
      17'd62918: data = 8'h02;
      17'd62919: data = 8'h04;
      17'd62920: data = 8'h05;
      17'd62921: data = 8'h05;
      17'd62922: data = 8'h02;
      17'd62923: data = 8'h02;
      17'd62924: data = 8'h01;
      17'd62925: data = 8'hfc;
      17'd62926: data = 8'hfd;
      17'd62927: data = 8'hfe;
      17'd62928: data = 8'hfd;
      17'd62929: data = 8'hfd;
      17'd62930: data = 8'h00;
      17'd62931: data = 8'h02;
      17'd62932: data = 8'h01;
      17'd62933: data = 8'hfe;
      17'd62934: data = 8'hfe;
      17'd62935: data = 8'hfd;
      17'd62936: data = 8'hf9;
      17'd62937: data = 8'hf6;
      17'd62938: data = 8'hf5;
      17'd62939: data = 8'hf9;
      17'd62940: data = 8'hf6;
      17'd62941: data = 8'hf5;
      17'd62942: data = 8'hf6;
      17'd62943: data = 8'hf6;
      17'd62944: data = 8'hf4;
      17'd62945: data = 8'hf1;
      17'd62946: data = 8'hf4;
      17'd62947: data = 8'hf1;
      17'd62948: data = 8'hef;
      17'd62949: data = 8'hf2;
      17'd62950: data = 8'hf5;
      17'd62951: data = 8'hf4;
      17'd62952: data = 8'hf4;
      17'd62953: data = 8'hf4;
      17'd62954: data = 8'hf5;
      17'd62955: data = 8'hf4;
      17'd62956: data = 8'hf2;
      17'd62957: data = 8'hf1;
      17'd62958: data = 8'hf1;
      17'd62959: data = 8'hf1;
      17'd62960: data = 8'hed;
      17'd62961: data = 8'hf4;
      17'd62962: data = 8'hf6;
      17'd62963: data = 8'hf5;
      17'd62964: data = 8'hf9;
      17'd62965: data = 8'hf5;
      17'd62966: data = 8'hf2;
      17'd62967: data = 8'hf1;
      17'd62968: data = 8'hf2;
      17'd62969: data = 8'hf5;
      17'd62970: data = 8'hf5;
      17'd62971: data = 8'hf5;
      17'd62972: data = 8'hf5;
      17'd62973: data = 8'hf9;
      17'd62974: data = 8'hfc;
      17'd62975: data = 8'hfa;
      17'd62976: data = 8'hf9;
      17'd62977: data = 8'hfc;
      17'd62978: data = 8'hfe;
      17'd62979: data = 8'h01;
      17'd62980: data = 8'h01;
      17'd62981: data = 8'h04;
      17'd62982: data = 8'h06;
      17'd62983: data = 8'h04;
      17'd62984: data = 8'h05;
      17'd62985: data = 8'h06;
      17'd62986: data = 8'h09;
      17'd62987: data = 8'h02;
      17'd62988: data = 8'h04;
      17'd62989: data = 8'h09;
      17'd62990: data = 8'h09;
      17'd62991: data = 8'h09;
      17'd62992: data = 8'h09;
      17'd62993: data = 8'h0d;
      17'd62994: data = 8'h12;
      17'd62995: data = 8'h13;
      17'd62996: data = 8'h0d;
      17'd62997: data = 8'h09;
      17'd62998: data = 8'h0c;
      17'd62999: data = 8'h0e;
      17'd63000: data = 8'h12;
      17'd63001: data = 8'h15;
      17'd63002: data = 8'h11;
      17'd63003: data = 8'h11;
      17'd63004: data = 8'h13;
      17'd63005: data = 8'h1a;
      17'd63006: data = 8'h19;
      17'd63007: data = 8'h13;
      17'd63008: data = 8'h13;
      17'd63009: data = 8'h16;
      17'd63010: data = 8'h1a;
      17'd63011: data = 8'h16;
      17'd63012: data = 8'h13;
      17'd63013: data = 8'h13;
      17'd63014: data = 8'h15;
      17'd63015: data = 8'h16;
      17'd63016: data = 8'h16;
      17'd63017: data = 8'h13;
      17'd63018: data = 8'h11;
      17'd63019: data = 8'h13;
      17'd63020: data = 8'h16;
      17'd63021: data = 8'h15;
      17'd63022: data = 8'h11;
      17'd63023: data = 8'h11;
      17'd63024: data = 8'h12;
      17'd63025: data = 8'h16;
      17'd63026: data = 8'h13;
      17'd63027: data = 8'h0e;
      17'd63028: data = 8'h11;
      17'd63029: data = 8'h11;
      17'd63030: data = 8'h11;
      17'd63031: data = 8'h0e;
      17'd63032: data = 8'h11;
      17'd63033: data = 8'h0e;
      17'd63034: data = 8'h0d;
      17'd63035: data = 8'h0d;
      17'd63036: data = 8'h0d;
      17'd63037: data = 8'h0d;
      17'd63038: data = 8'h0c;
      17'd63039: data = 8'h09;
      17'd63040: data = 8'h06;
      17'd63041: data = 8'h09;
      17'd63042: data = 8'h06;
      17'd63043: data = 8'h06;
      17'd63044: data = 8'h05;
      17'd63045: data = 8'h06;
      17'd63046: data = 8'h05;
      17'd63047: data = 8'h05;
      17'd63048: data = 8'h05;
      17'd63049: data = 8'h05;
      17'd63050: data = 8'h05;
      17'd63051: data = 8'h05;
      17'd63052: data = 8'h06;
      17'd63053: data = 8'h05;
      17'd63054: data = 8'h05;
      17'd63055: data = 8'h05;
      17'd63056: data = 8'h04;
      17'd63057: data = 8'h04;
      17'd63058: data = 8'h02;
      17'd63059: data = 8'h02;
      17'd63060: data = 8'h02;
      17'd63061: data = 8'hfe;
      17'd63062: data = 8'h00;
      17'd63063: data = 8'h00;
      17'd63064: data = 8'h00;
      17'd63065: data = 8'hfc;
      17'd63066: data = 8'hfc;
      17'd63067: data = 8'hfe;
      17'd63068: data = 8'hfd;
      17'd63069: data = 8'hfa;
      17'd63070: data = 8'hfc;
      17'd63071: data = 8'hfd;
      17'd63072: data = 8'hfd;
      17'd63073: data = 8'hfd;
      17'd63074: data = 8'hfe;
      17'd63075: data = 8'h01;
      17'd63076: data = 8'h00;
      17'd63077: data = 8'h00;
      17'd63078: data = 8'h01;
      17'd63079: data = 8'h01;
      17'd63080: data = 8'hfe;
      17'd63081: data = 8'hfc;
      17'd63082: data = 8'hfe;
      17'd63083: data = 8'hfe;
      17'd63084: data = 8'hfa;
      17'd63085: data = 8'hfa;
      17'd63086: data = 8'hfe;
      17'd63087: data = 8'h00;
      17'd63088: data = 8'hfd;
      17'd63089: data = 8'hfd;
      17'd63090: data = 8'h02;
      17'd63091: data = 8'h02;
      17'd63092: data = 8'h00;
      17'd63093: data = 8'hfe;
      17'd63094: data = 8'h01;
      17'd63095: data = 8'h00;
      17'd63096: data = 8'hfd;
      17'd63097: data = 8'hfe;
      17'd63098: data = 8'h00;
      17'd63099: data = 8'hfd;
      17'd63100: data = 8'hfc;
      17'd63101: data = 8'hfe;
      17'd63102: data = 8'hfe;
      17'd63103: data = 8'hfe;
      17'd63104: data = 8'hfd;
      17'd63105: data = 8'hfd;
      17'd63106: data = 8'hfd;
      17'd63107: data = 8'hf9;
      17'd63108: data = 8'hf6;
      17'd63109: data = 8'hfa;
      17'd63110: data = 8'hf6;
      17'd63111: data = 8'hf1;
      17'd63112: data = 8'hf1;
      17'd63113: data = 8'hf4;
      17'd63114: data = 8'hef;
      17'd63115: data = 8'hec;
      17'd63116: data = 8'hec;
      17'd63117: data = 8'hed;
      17'd63118: data = 8'hec;
      17'd63119: data = 8'hec;
      17'd63120: data = 8'hed;
      17'd63121: data = 8'hef;
      17'd63122: data = 8'hed;
      17'd63123: data = 8'hed;
      17'd63124: data = 8'hed;
      17'd63125: data = 8'hed;
      17'd63126: data = 8'hec;
      17'd63127: data = 8'he9;
      17'd63128: data = 8'heb;
      17'd63129: data = 8'heb;
      17'd63130: data = 8'he9;
      17'd63131: data = 8'he7;
      17'd63132: data = 8'heb;
      17'd63133: data = 8'heb;
      17'd63134: data = 8'heb;
      17'd63135: data = 8'heb;
      17'd63136: data = 8'heb;
      17'd63137: data = 8'heb;
      17'd63138: data = 8'heb;
      17'd63139: data = 8'hec;
      17'd63140: data = 8'hec;
      17'd63141: data = 8'hed;
      17'd63142: data = 8'hed;
      17'd63143: data = 8'hef;
      17'd63144: data = 8'hf2;
      17'd63145: data = 8'hf5;
      17'd63146: data = 8'hf6;
      17'd63147: data = 8'hf9;
      17'd63148: data = 8'hf6;
      17'd63149: data = 8'hf6;
      17'd63150: data = 8'hfa;
      17'd63151: data = 8'hfc;
      17'd63152: data = 8'hfa;
      17'd63153: data = 8'hfc;
      17'd63154: data = 8'hfc;
      17'd63155: data = 8'hfd;
      17'd63156: data = 8'hfd;
      17'd63157: data = 8'hfd;
      17'd63158: data = 8'hfd;
      17'd63159: data = 8'hfe;
      17'd63160: data = 8'h00;
      17'd63161: data = 8'hfe;
      17'd63162: data = 8'hfe;
      17'd63163: data = 8'h00;
      17'd63164: data = 8'h01;
      17'd63165: data = 8'h02;
      17'd63166: data = 8'h02;
      17'd63167: data = 8'h01;
      17'd63168: data = 8'h01;
      17'd63169: data = 8'h01;
      17'd63170: data = 8'h01;
      17'd63171: data = 8'h02;
      17'd63172: data = 8'h02;
      17'd63173: data = 8'h04;
      17'd63174: data = 8'h02;
      17'd63175: data = 8'h02;
      17'd63176: data = 8'h02;
      17'd63177: data = 8'h02;
      17'd63178: data = 8'h02;
      17'd63179: data = 8'h02;
      17'd63180: data = 8'h01;
      17'd63181: data = 8'h01;
      17'd63182: data = 8'h01;
      17'd63183: data = 8'h00;
      17'd63184: data = 8'h00;
      17'd63185: data = 8'h00;
      17'd63186: data = 8'h00;
      17'd63187: data = 8'h00;
      17'd63188: data = 8'h00;
      17'd63189: data = 8'hfe;
      17'd63190: data = 8'hfe;
      17'd63191: data = 8'hfe;
      17'd63192: data = 8'hfc;
      17'd63193: data = 8'hfd;
      17'd63194: data = 8'h00;
      17'd63195: data = 8'h00;
      17'd63196: data = 8'hfe;
      17'd63197: data = 8'hfe;
      17'd63198: data = 8'hfc;
      17'd63199: data = 8'hfc;
      17'd63200: data = 8'hfa;
      17'd63201: data = 8'hfa;
      17'd63202: data = 8'hf9;
      17'd63203: data = 8'hf6;
      17'd63204: data = 8'hfa;
      17'd63205: data = 8'hf6;
      17'd63206: data = 8'hf6;
      17'd63207: data = 8'hf5;
      17'd63208: data = 8'hf5;
      17'd63209: data = 8'hf6;
      17'd63210: data = 8'hf5;
      17'd63211: data = 8'hf5;
      17'd63212: data = 8'hf6;
      17'd63213: data = 8'hf5;
      17'd63214: data = 8'hf4;
      17'd63215: data = 8'hf4;
      17'd63216: data = 8'hf4;
      17'd63217: data = 8'hf9;
      17'd63218: data = 8'hf9;
      17'd63219: data = 8'hf6;
      17'd63220: data = 8'hf6;
      17'd63221: data = 8'hf6;
      17'd63222: data = 8'hf6;
      17'd63223: data = 8'hf6;
      17'd63224: data = 8'hf5;
      17'd63225: data = 8'hf4;
      17'd63226: data = 8'hf5;
      17'd63227: data = 8'hf5;
      17'd63228: data = 8'hf4;
      17'd63229: data = 8'hf2;
      17'd63230: data = 8'hf6;
      17'd63231: data = 8'hf6;
      17'd63232: data = 8'hfa;
      17'd63233: data = 8'hfa;
      17'd63234: data = 8'hf6;
      17'd63235: data = 8'hf9;
      17'd63236: data = 8'hfa;
      17'd63237: data = 8'hfc;
      17'd63238: data = 8'hfd;
      17'd63239: data = 8'hfc;
      17'd63240: data = 8'hfd;
      17'd63241: data = 8'h01;
      17'd63242: data = 8'h01;
      17'd63243: data = 8'h00;
      17'd63244: data = 8'h00;
      17'd63245: data = 8'h04;
      17'd63246: data = 8'h04;
      17'd63247: data = 8'h02;
      17'd63248: data = 8'h05;
      17'd63249: data = 8'h0a;
      17'd63250: data = 8'h06;
      17'd63251: data = 8'h02;
      17'd63252: data = 8'h05;
      17'd63253: data = 8'h0c;
      17'd63254: data = 8'h0a;
      17'd63255: data = 8'h06;
      17'd63256: data = 8'h06;
      17'd63257: data = 8'h0a;
      17'd63258: data = 8'h0e;
      17'd63259: data = 8'h11;
      17'd63260: data = 8'h0e;
      17'd63261: data = 8'h0e;
      17'd63262: data = 8'h12;
      17'd63263: data = 8'h15;
      17'd63264: data = 8'h16;
      17'd63265: data = 8'h13;
      17'd63266: data = 8'h11;
      17'd63267: data = 8'h12;
      17'd63268: data = 8'h19;
      17'd63269: data = 8'h1a;
      17'd63270: data = 8'h13;
      17'd63271: data = 8'h12;
      17'd63272: data = 8'h16;
      17'd63273: data = 8'h19;
      17'd63274: data = 8'h13;
      17'd63275: data = 8'h13;
      17'd63276: data = 8'h15;
      17'd63277: data = 8'h15;
      17'd63278: data = 8'h13;
      17'd63279: data = 8'h15;
      17'd63280: data = 8'h15;
      17'd63281: data = 8'h16;
      17'd63282: data = 8'h13;
      17'd63283: data = 8'h12;
      17'd63284: data = 8'h15;
      17'd63285: data = 8'h16;
      17'd63286: data = 8'h11;
      17'd63287: data = 8'h0e;
      17'd63288: data = 8'h13;
      17'd63289: data = 8'h13;
      17'd63290: data = 8'h13;
      17'd63291: data = 8'h0e;
      17'd63292: data = 8'h0d;
      17'd63293: data = 8'h0d;
      17'd63294: data = 8'h0e;
      17'd63295: data = 8'h11;
      17'd63296: data = 8'h0d;
      17'd63297: data = 8'h0c;
      17'd63298: data = 8'h0a;
      17'd63299: data = 8'h0a;
      17'd63300: data = 8'h0a;
      17'd63301: data = 8'h06;
      17'd63302: data = 8'h06;
      17'd63303: data = 8'h05;
      17'd63304: data = 8'h06;
      17'd63305: data = 8'h06;
      17'd63306: data = 8'h06;
      17'd63307: data = 8'h06;
      17'd63308: data = 8'h06;
      17'd63309: data = 8'h06;
      17'd63310: data = 8'h05;
      17'd63311: data = 8'h09;
      17'd63312: data = 8'h05;
      17'd63313: data = 8'h04;
      17'd63314: data = 8'h01;
      17'd63315: data = 8'h01;
      17'd63316: data = 8'h00;
      17'd63317: data = 8'h00;
      17'd63318: data = 8'h02;
      17'd63319: data = 8'hfe;
      17'd63320: data = 8'hfd;
      17'd63321: data = 8'h00;
      17'd63322: data = 8'h00;
      17'd63323: data = 8'hfe;
      17'd63324: data = 8'hfa;
      17'd63325: data = 8'hfd;
      17'd63326: data = 8'h01;
      17'd63327: data = 8'hfe;
      17'd63328: data = 8'hfc;
      17'd63329: data = 8'hfd;
      17'd63330: data = 8'hfd;
      17'd63331: data = 8'hfd;
      17'd63332: data = 8'hfe;
      17'd63333: data = 8'hfc;
      17'd63334: data = 8'hfc;
      17'd63335: data = 8'hfa;
      17'd63336: data = 8'hfc;
      17'd63337: data = 8'hfd;
      17'd63338: data = 8'hfa;
      17'd63339: data = 8'hf9;
      17'd63340: data = 8'hf9;
      17'd63341: data = 8'hfc;
      17'd63342: data = 8'hfa;
      17'd63343: data = 8'hf9;
      17'd63344: data = 8'hf9;
      17'd63345: data = 8'hf9;
      17'd63346: data = 8'hf5;
      17'd63347: data = 8'hf5;
      17'd63348: data = 8'hf6;
      17'd63349: data = 8'hf6;
      17'd63350: data = 8'hf4;
      17'd63351: data = 8'hf5;
      17'd63352: data = 8'hf5;
      17'd63353: data = 8'hf9;
      17'd63354: data = 8'hf6;
      17'd63355: data = 8'hf5;
      17'd63356: data = 8'hf5;
      17'd63357: data = 8'hf6;
      17'd63358: data = 8'hf9;
      17'd63359: data = 8'hf6;
      17'd63360: data = 8'hf6;
      17'd63361: data = 8'hf6;
      17'd63362: data = 8'hf6;
      17'd63363: data = 8'hfa;
      17'd63364: data = 8'hf6;
      17'd63365: data = 8'hf5;
      17'd63366: data = 8'hf9;
      17'd63367: data = 8'hfa;
      17'd63368: data = 8'hf9;
      17'd63369: data = 8'hf9;
      17'd63370: data = 8'hf9;
      17'd63371: data = 8'hf9;
      17'd63372: data = 8'hf9;
      17'd63373: data = 8'hf6;
      17'd63374: data = 8'hf9;
      17'd63375: data = 8'hfa;
      17'd63376: data = 8'hf9;
      17'd63377: data = 8'hf9;
      17'd63378: data = 8'hf9;
      17'd63379: data = 8'hfa;
      17'd63380: data = 8'hf9;
      17'd63381: data = 8'hfa;
      17'd63382: data = 8'hf9;
      17'd63383: data = 8'hf9;
      17'd63384: data = 8'hf6;
      17'd63385: data = 8'hf6;
      17'd63386: data = 8'hf6;
      17'd63387: data = 8'hf5;
      17'd63388: data = 8'hf4;
      17'd63389: data = 8'hf4;
      17'd63390: data = 8'hf2;
      17'd63391: data = 8'hef;
      17'd63392: data = 8'hf1;
      17'd63393: data = 8'hf1;
      17'd63394: data = 8'hef;
      17'd63395: data = 8'hf1;
      17'd63396: data = 8'hed;
      17'd63397: data = 8'hed;
      17'd63398: data = 8'hec;
      17'd63399: data = 8'hed;
      17'd63400: data = 8'hec;
      17'd63401: data = 8'hec;
      17'd63402: data = 8'hec;
      17'd63403: data = 8'hec;
      17'd63404: data = 8'hec;
      17'd63405: data = 8'heb;
      17'd63406: data = 8'hec;
      17'd63407: data = 8'hec;
      17'd63408: data = 8'hec;
      17'd63409: data = 8'hef;
      17'd63410: data = 8'hef;
      17'd63411: data = 8'hef;
      17'd63412: data = 8'hf1;
      17'd63413: data = 8'hef;
      17'd63414: data = 8'hef;
      17'd63415: data = 8'hef;
      17'd63416: data = 8'hf1;
      17'd63417: data = 8'hef;
      17'd63418: data = 8'hef;
      17'd63419: data = 8'hf2;
      17'd63420: data = 8'hf2;
      17'd63421: data = 8'hf4;
      17'd63422: data = 8'hf5;
      17'd63423: data = 8'hf6;
      17'd63424: data = 8'hf9;
      17'd63425: data = 8'hfa;
      17'd63426: data = 8'hfa;
      17'd63427: data = 8'hfa;
      17'd63428: data = 8'hfc;
      17'd63429: data = 8'hf9;
      17'd63430: data = 8'hfc;
      17'd63431: data = 8'hfc;
      17'd63432: data = 8'hfd;
      17'd63433: data = 8'hfd;
      17'd63434: data = 8'hfe;
      17'd63435: data = 8'h00;
      17'd63436: data = 8'h01;
      17'd63437: data = 8'h02;
      17'd63438: data = 8'h02;
      17'd63439: data = 8'h04;
      17'd63440: data = 8'h05;
      17'd63441: data = 8'h05;
      17'd63442: data = 8'h05;
      17'd63443: data = 8'h05;
      17'd63444: data = 8'h04;
      17'd63445: data = 8'h01;
      17'd63446: data = 8'h01;
      17'd63447: data = 8'h04;
      17'd63448: data = 8'h02;
      17'd63449: data = 8'h01;
      17'd63450: data = 8'h04;
      17'd63451: data = 8'h05;
      17'd63452: data = 8'h05;
      17'd63453: data = 8'h04;
      17'd63454: data = 8'h05;
      17'd63455: data = 8'h06;
      17'd63456: data = 8'h09;
      17'd63457: data = 8'h05;
      17'd63458: data = 8'h09;
      17'd63459: data = 8'h06;
      17'd63460: data = 8'h06;
      17'd63461: data = 8'h06;
      17'd63462: data = 8'h05;
      17'd63463: data = 8'h06;
      17'd63464: data = 8'h05;
      17'd63465: data = 8'h05;
      17'd63466: data = 8'h05;
      17'd63467: data = 8'h09;
      17'd63468: data = 8'h05;
      17'd63469: data = 8'h06;
      17'd63470: data = 8'h09;
      17'd63471: data = 8'h09;
      17'd63472: data = 8'h06;
      17'd63473: data = 8'h05;
      17'd63474: data = 8'h04;
      17'd63475: data = 8'h02;
      17'd63476: data = 8'h01;
      17'd63477: data = 8'h04;
      17'd63478: data = 8'h04;
      17'd63479: data = 8'h02;
      17'd63480: data = 8'h02;
      17'd63481: data = 8'h02;
      17'd63482: data = 8'h06;
      17'd63483: data = 8'h04;
      17'd63484: data = 8'h05;
      17'd63485: data = 8'h06;
      17'd63486: data = 8'h05;
      17'd63487: data = 8'h05;
      17'd63488: data = 8'h05;
      17'd63489: data = 8'h06;
      17'd63490: data = 8'h05;
      17'd63491: data = 8'h02;
      17'd63492: data = 8'h01;
      17'd63493: data = 8'h02;
      17'd63494: data = 8'h01;
      17'd63495: data = 8'hfe;
      17'd63496: data = 8'h00;
      17'd63497: data = 8'h02;
      17'd63498: data = 8'h05;
      17'd63499: data = 8'h02;
      17'd63500: data = 8'h01;
      17'd63501: data = 8'h01;
      17'd63502: data = 8'h02;
      17'd63503: data = 8'h00;
      17'd63504: data = 8'hfd;
      17'd63505: data = 8'hfc;
      17'd63506: data = 8'hfe;
      17'd63507: data = 8'h00;
      17'd63508: data = 8'h00;
      17'd63509: data = 8'hfe;
      17'd63510: data = 8'hfd;
      17'd63511: data = 8'h02;
      17'd63512: data = 8'h04;
      17'd63513: data = 8'h04;
      17'd63514: data = 8'hfe;
      17'd63515: data = 8'hfd;
      17'd63516: data = 8'h02;
      17'd63517: data = 8'h01;
      17'd63518: data = 8'hfe;
      17'd63519: data = 8'hfa;
      17'd63520: data = 8'hfc;
      17'd63521: data = 8'h00;
      17'd63522: data = 8'h01;
      17'd63523: data = 8'hfe;
      17'd63524: data = 8'hfd;
      17'd63525: data = 8'h00;
      17'd63526: data = 8'h04;
      17'd63527: data = 8'h05;
      17'd63528: data = 8'h02;
      17'd63529: data = 8'h01;
      17'd63530: data = 8'h05;
      17'd63531: data = 8'h06;
      17'd63532: data = 8'h06;
      17'd63533: data = 8'h05;
      17'd63534: data = 8'h05;
      17'd63535: data = 8'h04;
      17'd63536: data = 8'h04;
      17'd63537: data = 8'h09;
      17'd63538: data = 8'h06;
      17'd63539: data = 8'h05;
      17'd63540: data = 8'h06;
      17'd63541: data = 8'h0c;
      17'd63542: data = 8'h11;
      17'd63543: data = 8'h0e;
      17'd63544: data = 8'h0c;
      17'd63545: data = 8'h0d;
      17'd63546: data = 8'h0e;
      17'd63547: data = 8'h0e;
      17'd63548: data = 8'h11;
      17'd63549: data = 8'h12;
      17'd63550: data = 8'h11;
      17'd63551: data = 8'h11;
      17'd63552: data = 8'h12;
      17'd63553: data = 8'h13;
      17'd63554: data = 8'h11;
      17'd63555: data = 8'h0d;
      17'd63556: data = 8'h0e;
      17'd63557: data = 8'h12;
      17'd63558: data = 8'h12;
      17'd63559: data = 8'h12;
      17'd63560: data = 8'h11;
      17'd63561: data = 8'h12;
      17'd63562: data = 8'h11;
      17'd63563: data = 8'h0e;
      17'd63564: data = 8'h11;
      17'd63565: data = 8'h0e;
      17'd63566: data = 8'h0e;
      17'd63567: data = 8'h11;
      17'd63568: data = 8'h0e;
      17'd63569: data = 8'h0d;
      17'd63570: data = 8'h0d;
      17'd63571: data = 8'h0d;
      17'd63572: data = 8'h0d;
      17'd63573: data = 8'h0a;
      17'd63574: data = 8'h0a;
      17'd63575: data = 8'h0c;
      17'd63576: data = 8'h09;
      17'd63577: data = 8'h05;
      17'd63578: data = 8'h05;
      17'd63579: data = 8'h06;
      17'd63580: data = 8'h06;
      17'd63581: data = 8'h04;
      17'd63582: data = 8'h02;
      17'd63583: data = 8'h04;
      17'd63584: data = 8'h02;
      17'd63585: data = 8'h01;
      17'd63586: data = 8'h02;
      17'd63587: data = 8'h02;
      17'd63588: data = 8'h00;
      17'd63589: data = 8'hfe;
      17'd63590: data = 8'hfe;
      17'd63591: data = 8'hfe;
      17'd63592: data = 8'hfe;
      17'd63593: data = 8'h00;
      17'd63594: data = 8'h00;
      17'd63595: data = 8'hfc;
      17'd63596: data = 8'hfa;
      17'd63597: data = 8'hf9;
      17'd63598: data = 8'hfa;
      17'd63599: data = 8'hf6;
      17'd63600: data = 8'hf9;
      17'd63601: data = 8'hfc;
      17'd63602: data = 8'hf9;
      17'd63603: data = 8'hf9;
      17'd63604: data = 8'hf6;
      17'd63605: data = 8'hf6;
      17'd63606: data = 8'hf9;
      17'd63607: data = 8'hf6;
      17'd63608: data = 8'hf5;
      17'd63609: data = 8'hf6;
      17'd63610: data = 8'hf9;
      17'd63611: data = 8'hf5;
      17'd63612: data = 8'hf4;
      17'd63613: data = 8'hf5;
      17'd63614: data = 8'hf6;
      17'd63615: data = 8'hf4;
      17'd63616: data = 8'hf2;
      17'd63617: data = 8'hf2;
      17'd63618: data = 8'hf2;
      17'd63619: data = 8'hf2;
      17'd63620: data = 8'hf4;
      17'd63621: data = 8'hf2;
      17'd63622: data = 8'hf2;
      17'd63623: data = 8'hf4;
      17'd63624: data = 8'hf2;
      17'd63625: data = 8'hf1;
      17'd63626: data = 8'hef;
      17'd63627: data = 8'hef;
      17'd63628: data = 8'hef;
      17'd63629: data = 8'hed;
      17'd63630: data = 8'hef;
      17'd63631: data = 8'hef;
      17'd63632: data = 8'hef;
      17'd63633: data = 8'hef;
      17'd63634: data = 8'hf1;
      17'd63635: data = 8'hf2;
      17'd63636: data = 8'hf2;
      17'd63637: data = 8'hf2;
      17'd63638: data = 8'hf2;
      17'd63639: data = 8'hf1;
      17'd63640: data = 8'hf1;
      17'd63641: data = 8'hf2;
      17'd63642: data = 8'hf1;
      17'd63643: data = 8'hf2;
      17'd63644: data = 8'hf2;
      17'd63645: data = 8'hf2;
      17'd63646: data = 8'hf4;
      17'd63647: data = 8'hf4;
      17'd63648: data = 8'hf4;
      17'd63649: data = 8'hf4;
      17'd63650: data = 8'hf5;
      17'd63651: data = 8'hf9;
      17'd63652: data = 8'hfa;
      17'd63653: data = 8'hf6;
      17'd63654: data = 8'hfa;
      17'd63655: data = 8'hf9;
      17'd63656: data = 8'hf9;
      17'd63657: data = 8'hf6;
      17'd63658: data = 8'hf6;
      17'd63659: data = 8'hf9;
      17'd63660: data = 8'hf9;
      17'd63661: data = 8'hf9;
      17'd63662: data = 8'hfa;
      17'd63663: data = 8'hfc;
      17'd63664: data = 8'hfe;
      17'd63665: data = 8'h00;
      17'd63666: data = 8'h00;
      17'd63667: data = 8'h00;
      17'd63668: data = 8'h00;
      17'd63669: data = 8'hfd;
      17'd63670: data = 8'hfc;
      17'd63671: data = 8'hfd;
      17'd63672: data = 8'hfd;
      17'd63673: data = 8'hfd;
      17'd63674: data = 8'hfd;
      17'd63675: data = 8'hfd;
      17'd63676: data = 8'hfe;
      17'd63677: data = 8'h00;
      17'd63678: data = 8'hfd;
      17'd63679: data = 8'hfd;
      17'd63680: data = 8'hfd;
      17'd63681: data = 8'hfd;
      17'd63682: data = 8'hfe;
      17'd63683: data = 8'hfd;
      17'd63684: data = 8'hfd;
      17'd63685: data = 8'hfc;
      17'd63686: data = 8'hfa;
      17'd63687: data = 8'hfc;
      17'd63688: data = 8'hfa;
      17'd63689: data = 8'hfa;
      17'd63690: data = 8'hf9;
      17'd63691: data = 8'hf9;
      17'd63692: data = 8'hfa;
      17'd63693: data = 8'hfa;
      17'd63694: data = 8'hfa;
      17'd63695: data = 8'hf9;
      17'd63696: data = 8'hf9;
      17'd63697: data = 8'hfa;
      17'd63698: data = 8'hfc;
      17'd63699: data = 8'hf9;
      17'd63700: data = 8'hf6;
      17'd63701: data = 8'hf6;
      17'd63702: data = 8'hf9;
      17'd63703: data = 8'hfa;
      17'd63704: data = 8'hfa;
      17'd63705: data = 8'hf5;
      17'd63706: data = 8'hf9;
      17'd63707: data = 8'hfc;
      17'd63708: data = 8'hfc;
      17'd63709: data = 8'hfd;
      17'd63710: data = 8'hfd;
      17'd63711: data = 8'hfc;
      17'd63712: data = 8'hfd;
      17'd63713: data = 8'hfd;
      17'd63714: data = 8'hfd;
      17'd63715: data = 8'hfe;
      17'd63716: data = 8'hfc;
      17'd63717: data = 8'hfd;
      17'd63718: data = 8'hfd;
      17'd63719: data = 8'hfc;
      17'd63720: data = 8'hfc;
      17'd63721: data = 8'hfd;
      17'd63722: data = 8'hfd;
      17'd63723: data = 8'hfe;
      17'd63724: data = 8'h00;
      17'd63725: data = 8'h00;
      17'd63726: data = 8'h01;
      17'd63727: data = 8'h00;
      17'd63728: data = 8'h00;
      17'd63729: data = 8'h01;
      17'd63730: data = 8'h00;
      17'd63731: data = 8'h01;
      17'd63732: data = 8'h02;
      17'd63733: data = 8'h02;
      17'd63734: data = 8'h04;
      17'd63735: data = 8'h02;
      17'd63736: data = 8'h01;
      17'd63737: data = 8'h02;
      17'd63738: data = 8'h05;
      17'd63739: data = 8'h04;
      17'd63740: data = 8'h04;
      17'd63741: data = 8'h02;
      17'd63742: data = 8'h04;
      17'd63743: data = 8'h02;
      17'd63744: data = 8'h02;
      17'd63745: data = 8'h05;
      17'd63746: data = 8'h04;
      17'd63747: data = 8'h05;
      17'd63748: data = 8'h04;
      17'd63749: data = 8'h04;
      17'd63750: data = 8'h05;
      17'd63751: data = 8'h04;
      17'd63752: data = 8'h04;
      17'd63753: data = 8'h06;
      17'd63754: data = 8'h06;
      17'd63755: data = 8'h06;
      17'd63756: data = 8'h06;
      17'd63757: data = 8'h05;
      17'd63758: data = 8'h06;
      17'd63759: data = 8'h09;
      17'd63760: data = 8'h09;
      17'd63761: data = 8'h09;
      17'd63762: data = 8'h09;
      17'd63763: data = 8'h05;
      17'd63764: data = 8'h05;
      17'd63765: data = 8'h05;
      17'd63766: data = 8'h05;
      17'd63767: data = 8'h05;
      17'd63768: data = 8'h06;
      17'd63769: data = 8'h05;
      17'd63770: data = 8'h06;
      17'd63771: data = 8'h09;
      17'd63772: data = 8'h06;
      17'd63773: data = 8'h05;
      17'd63774: data = 8'h06;
      17'd63775: data = 8'h05;
      17'd63776: data = 8'h05;
      17'd63777: data = 8'h05;
      17'd63778: data = 8'h05;
      17'd63779: data = 8'h05;
      17'd63780: data = 8'h04;
      17'd63781: data = 8'h04;
      17'd63782: data = 8'h05;
      17'd63783: data = 8'h06;
      17'd63784: data = 8'h05;
      17'd63785: data = 8'h05;
      17'd63786: data = 8'h09;
      17'd63787: data = 8'h06;
      17'd63788: data = 8'h06;
      17'd63789: data = 8'h06;
      17'd63790: data = 8'h05;
      17'd63791: data = 8'h05;
      17'd63792: data = 8'h05;
      17'd63793: data = 8'h04;
      17'd63794: data = 8'h01;
      17'd63795: data = 8'h00;
      17'd63796: data = 8'h01;
      17'd63797: data = 8'h01;
      17'd63798: data = 8'h00;
      17'd63799: data = 8'h00;
      17'd63800: data = 8'h01;
      17'd63801: data = 8'h02;
      17'd63802: data = 8'h02;
      17'd63803: data = 8'h02;
      17'd63804: data = 8'h01;
      17'd63805: data = 8'h02;
      17'd63806: data = 8'h02;
      17'd63807: data = 8'h01;
      17'd63808: data = 8'h01;
      17'd63809: data = 8'h00;
      17'd63810: data = 8'hfe;
      17'd63811: data = 8'hfe;
      17'd63812: data = 8'hfe;
      17'd63813: data = 8'hfe;
      17'd63814: data = 8'hfe;
      17'd63815: data = 8'hfe;
      17'd63816: data = 8'hfe;
      17'd63817: data = 8'hfe;
      17'd63818: data = 8'h00;
      17'd63819: data = 8'h00;
      17'd63820: data = 8'hfe;
      17'd63821: data = 8'h00;
      17'd63822: data = 8'h00;
      17'd63823: data = 8'hfe;
      17'd63824: data = 8'h00;
      17'd63825: data = 8'h00;
      17'd63826: data = 8'h00;
      17'd63827: data = 8'hfe;
      17'd63828: data = 8'hfd;
      17'd63829: data = 8'hfd;
      17'd63830: data = 8'hfe;
      17'd63831: data = 8'h00;
      17'd63832: data = 8'h01;
      17'd63833: data = 8'h01;
      17'd63834: data = 8'h02;
      17'd63835: data = 8'h04;
      17'd63836: data = 8'h02;
      17'd63837: data = 8'h02;
      17'd63838: data = 8'h00;
      17'd63839: data = 8'h00;
      17'd63840: data = 8'h01;
      17'd63841: data = 8'h00;
      17'd63842: data = 8'h00;
      17'd63843: data = 8'h01;
      17'd63844: data = 8'h00;
      17'd63845: data = 8'h01;
      17'd63846: data = 8'h02;
      17'd63847: data = 8'h02;
      17'd63848: data = 8'h04;
      17'd63849: data = 8'h02;
      17'd63850: data = 8'h02;
      17'd63851: data = 8'h02;
      17'd63852: data = 8'h05;
      17'd63853: data = 8'h05;
      17'd63854: data = 8'h04;
      17'd63855: data = 8'h02;
      17'd63856: data = 8'h02;
      17'd63857: data = 8'h04;
      17'd63858: data = 8'h02;
      17'd63859: data = 8'h01;
      17'd63860: data = 8'h01;
      17'd63861: data = 8'h01;
      17'd63862: data = 8'h02;
      17'd63863: data = 8'h02;
      17'd63864: data = 8'h04;
      17'd63865: data = 8'h05;
      17'd63866: data = 8'h05;
      17'd63867: data = 8'h05;
      17'd63868: data = 8'h05;
      17'd63869: data = 8'h04;
      17'd63870: data = 8'h04;
      17'd63871: data = 8'h02;
      17'd63872: data = 8'h02;
      17'd63873: data = 8'h02;
      17'd63874: data = 8'h02;
      17'd63875: data = 8'h02;
      17'd63876: data = 8'h01;
      17'd63877: data = 8'h00;
      17'd63878: data = 8'h00;
      17'd63879: data = 8'h01;
      17'd63880: data = 8'hfe;
      17'd63881: data = 8'hfe;
      17'd63882: data = 8'h01;
      17'd63883: data = 8'h00;
      17'd63884: data = 8'h00;
      17'd63885: data = 8'h00;
      17'd63886: data = 8'h00;
      17'd63887: data = 8'hfe;
      17'd63888: data = 8'h00;
      17'd63889: data = 8'hfe;
      17'd63890: data = 8'h00;
      17'd63891: data = 8'hfe;
      17'd63892: data = 8'hfd;
      17'd63893: data = 8'hfc;
      17'd63894: data = 8'hfc;
      17'd63895: data = 8'hfe;
      17'd63896: data = 8'hfd;
      17'd63897: data = 8'hfa;
      17'd63898: data = 8'hfa;
      17'd63899: data = 8'hfc;
      17'd63900: data = 8'hfd;
      17'd63901: data = 8'hfd;
      17'd63902: data = 8'hfc;
      17'd63903: data = 8'hfa;
      17'd63904: data = 8'hfa;
      17'd63905: data = 8'hf9;
      17'd63906: data = 8'hf5;
      17'd63907: data = 8'hf6;
      17'd63908: data = 8'hf6;
      17'd63909: data = 8'hf9;
      17'd63910: data = 8'hfa;
      17'd63911: data = 8'hf6;
      17'd63912: data = 8'hf6;
      17'd63913: data = 8'hf6;
      17'd63914: data = 8'hf5;
      17'd63915: data = 8'hf6;
      17'd63916: data = 8'hf6;
      17'd63917: data = 8'hf9;
      17'd63918: data = 8'hf9;
      17'd63919: data = 8'hf6;
      17'd63920: data = 8'hf6;
      17'd63921: data = 8'hf6;
      17'd63922: data = 8'hf9;
      17'd63923: data = 8'hfa;
      17'd63924: data = 8'hf6;
      17'd63925: data = 8'hf6;
      17'd63926: data = 8'hfa;
      17'd63927: data = 8'hf9;
      17'd63928: data = 8'hfa;
      17'd63929: data = 8'hfc;
      17'd63930: data = 8'hfa;
      17'd63931: data = 8'hfc;
      17'd63932: data = 8'hfc;
      17'd63933: data = 8'hfc;
      17'd63934: data = 8'hfc;
      17'd63935: data = 8'hfc;
      17'd63936: data = 8'hfc;
      17'd63937: data = 8'hfc;
      17'd63938: data = 8'hfa;
      17'd63939: data = 8'hfa;
      17'd63940: data = 8'hfa;
      17'd63941: data = 8'hf9;
      17'd63942: data = 8'hfa;
      17'd63943: data = 8'hfd;
      17'd63944: data = 8'hfc;
      17'd63945: data = 8'hfa;
      17'd63946: data = 8'hfd;
      17'd63947: data = 8'hfc;
      17'd63948: data = 8'hfc;
      17'd63949: data = 8'hfa;
      17'd63950: data = 8'hfc;
      17'd63951: data = 8'hfd;
      17'd63952: data = 8'hfd;
      17'd63953: data = 8'hfd;
      17'd63954: data = 8'hfe;
      17'd63955: data = 8'hfc;
      17'd63956: data = 8'hfd;
      17'd63957: data = 8'hfc;
      17'd63958: data = 8'hfa;
      17'd63959: data = 8'hfc;
      17'd63960: data = 8'hfc;
      17'd63961: data = 8'hfc;
      17'd63962: data = 8'hfc;
      17'd63963: data = 8'hfc;
      17'd63964: data = 8'hfd;
      17'd63965: data = 8'hfe;
      17'd63966: data = 8'hfe;
      17'd63967: data = 8'hfd;
      17'd63968: data = 8'hfd;
      17'd63969: data = 8'hfd;
      17'd63970: data = 8'hfd;
      17'd63971: data = 8'hfe;
      17'd63972: data = 8'h00;
      17'd63973: data = 8'h00;
      17'd63974: data = 8'h00;
      17'd63975: data = 8'h00;
      17'd63976: data = 8'h00;
      17'd63977: data = 8'hfe;
      17'd63978: data = 8'hfe;
      17'd63979: data = 8'hfe;
      17'd63980: data = 8'hfe;
      17'd63981: data = 8'hfe;
      17'd63982: data = 8'hfd;
      17'd63983: data = 8'hfd;
      17'd63984: data = 8'hfd;
      17'd63985: data = 8'hfd;
      17'd63986: data = 8'hfe;
      17'd63987: data = 8'hfd;
      17'd63988: data = 8'hfd;
      17'd63989: data = 8'hfd;
      17'd63990: data = 8'hfe;
      17'd63991: data = 8'h00;
      17'd63992: data = 8'h01;
      17'd63993: data = 8'h02;
      17'd63994: data = 8'h01;
      17'd63995: data = 8'h00;
      17'd63996: data = 8'h00;
      17'd63997: data = 8'h00;
      17'd63998: data = 8'h00;
      17'd63999: data = 8'h00;
      17'd64000: data = 8'h00;
      17'd64001: data = 8'h00;
      17'd64002: data = 8'h01;
      17'd64003: data = 8'h00;
      17'd64004: data = 8'h00;
      17'd64005: data = 8'h02;
      17'd64006: data = 8'h00;
      17'd64007: data = 8'h01;
      17'd64008: data = 8'h02;
      17'd64009: data = 8'h01;
      17'd64010: data = 8'h02;
      17'd64011: data = 8'h02;
      17'd64012: data = 8'h02;
      17'd64013: data = 8'h01;
      17'd64014: data = 8'h02;
      17'd64015: data = 8'h01;
      17'd64016: data = 8'h01;
      17'd64017: data = 8'h01;
      17'd64018: data = 8'h01;
      17'd64019: data = 8'h01;
      17'd64020: data = 8'h04;
      17'd64021: data = 8'h04;
      17'd64022: data = 8'h01;
      17'd64023: data = 8'h02;
      17'd64024: data = 8'h02;
      17'd64025: data = 8'h01;
      17'd64026: data = 8'h02;
      17'd64027: data = 8'h02;
      17'd64028: data = 8'h01;
      17'd64029: data = 8'h04;
      17'd64030: data = 8'h02;
      17'd64031: data = 8'h01;
      17'd64032: data = 8'h01;
      17'd64033: data = 8'h02;
      17'd64034: data = 8'h02;
      17'd64035: data = 8'h02;
      17'd64036: data = 8'h01;
      17'd64037: data = 8'h02;
      17'd64038: data = 8'h04;
      17'd64039: data = 8'h02;
      17'd64040: data = 8'h02;
      17'd64041: data = 8'h02;
      17'd64042: data = 8'h04;
      17'd64043: data = 8'h04;
      17'd64044: data = 8'h04;
      17'd64045: data = 8'h04;
      17'd64046: data = 8'h02;
      17'd64047: data = 8'h04;
      17'd64048: data = 8'h02;
      17'd64049: data = 8'h01;
      17'd64050: data = 8'h02;
      17'd64051: data = 8'h01;
      17'd64052: data = 8'h02;
      17'd64053: data = 8'h01;
      17'd64054: data = 8'h04;
      17'd64055: data = 8'h04;
      17'd64056: data = 8'h04;
      17'd64057: data = 8'h06;
      17'd64058: data = 8'h02;
      17'd64059: data = 8'h05;
      17'd64060: data = 8'h05;
      17'd64061: data = 8'h02;
      17'd64062: data = 8'h02;
      17'd64063: data = 8'h02;
      17'd64064: data = 8'h02;
      17'd64065: data = 8'h01;
      17'd64066: data = 8'h02;
      17'd64067: data = 8'h04;
      17'd64068: data = 8'h02;
      17'd64069: data = 8'h01;
      17'd64070: data = 8'h02;
      17'd64071: data = 8'h01;
      17'd64072: data = 8'h02;
      17'd64073: data = 8'h04;
      17'd64074: data = 8'h04;
      17'd64075: data = 8'h04;
      17'd64076: data = 8'h01;
      17'd64077: data = 8'h02;
      17'd64078: data = 8'h02;
      17'd64079: data = 8'h00;
      17'd64080: data = 8'h01;
      17'd64081: data = 8'h02;
      17'd64082: data = 8'h01;
      17'd64083: data = 8'h01;
      17'd64084: data = 8'h02;
      17'd64085: data = 8'h01;
      17'd64086: data = 8'h01;
      17'd64087: data = 8'h02;
      17'd64088: data = 8'h02;
      17'd64089: data = 8'h02;
      17'd64090: data = 8'h01;
      17'd64091: data = 8'h01;
      17'd64092: data = 8'h01;
      17'd64093: data = 8'hfe;
      17'd64094: data = 8'hfe;
      17'd64095: data = 8'h00;
      17'd64096: data = 8'h02;
      17'd64097: data = 8'h01;
      17'd64098: data = 8'h01;
      17'd64099: data = 8'h02;
      17'd64100: data = 8'h02;
      17'd64101: data = 8'h01;
      17'd64102: data = 8'h01;
      17'd64103: data = 8'h02;
      17'd64104: data = 8'h01;
      17'd64105: data = 8'h01;
      17'd64106: data = 8'h02;
      17'd64107: data = 8'h02;
      17'd64108: data = 8'h02;
      17'd64109: data = 8'h02;
      17'd64110: data = 8'h01;
      17'd64111: data = 8'h02;
      17'd64112: data = 8'h01;
      17'd64113: data = 8'h00;
      17'd64114: data = 8'h00;
      17'd64115: data = 8'h00;
      17'd64116: data = 8'h04;
      17'd64117: data = 8'h01;
      17'd64118: data = 8'h04;
      17'd64119: data = 8'h01;
      17'd64120: data = 8'h01;
      17'd64121: data = 8'h01;
      17'd64122: data = 8'hfe;
      17'd64123: data = 8'h00;
      17'd64124: data = 8'hfe;
      17'd64125: data = 8'h00;
      17'd64126: data = 8'hfe;
      17'd64127: data = 8'hfe;
      17'd64128: data = 8'h00;
      17'd64129: data = 8'h01;
      17'd64130: data = 8'h00;
      17'd64131: data = 8'h00;
      17'd64132: data = 8'h00;
      17'd64133: data = 8'hfe;
      17'd64134: data = 8'hfe;
      17'd64135: data = 8'hfe;
      17'd64136: data = 8'hfe;
      17'd64137: data = 8'hfd;
      17'd64138: data = 8'hfe;
      17'd64139: data = 8'hfe;
      17'd64140: data = 8'hfd;
      17'd64141: data = 8'hfe;
      17'd64142: data = 8'hfe;
      17'd64143: data = 8'hfe;
      17'd64144: data = 8'h00;
      17'd64145: data = 8'h00;
      17'd64146: data = 8'hfd;
      17'd64147: data = 8'hfd;
      17'd64148: data = 8'hfe;
      17'd64149: data = 8'hfe;
      17'd64150: data = 8'hfe;
      17'd64151: data = 8'hfe;
      17'd64152: data = 8'hfe;
      17'd64153: data = 8'hfd;
      17'd64154: data = 8'hfe;
      17'd64155: data = 8'hfe;
      17'd64156: data = 8'hfe;
      17'd64157: data = 8'h01;
      17'd64158: data = 8'h00;
      17'd64159: data = 8'hfe;
      17'd64160: data = 8'h00;
      17'd64161: data = 8'h00;
      17'd64162: data = 8'h00;
      17'd64163: data = 8'h00;
      17'd64164: data = 8'hfe;
      17'd64165: data = 8'hfd;
      17'd64166: data = 8'hfd;
      17'd64167: data = 8'hfd;
      17'd64168: data = 8'hfe;
      17'd64169: data = 8'h01;
      17'd64170: data = 8'h01;
      17'd64171: data = 8'h01;
      17'd64172: data = 8'h00;
      17'd64173: data = 8'h01;
      17'd64174: data = 8'h01;
      17'd64175: data = 8'h00;
      17'd64176: data = 8'h00;
      17'd64177: data = 8'h00;
      17'd64178: data = 8'h01;
      17'd64179: data = 8'h01;
      17'd64180: data = 8'h00;
      17'd64181: data = 8'h00;
      17'd64182: data = 8'h00;
      17'd64183: data = 8'h00;
      17'd64184: data = 8'h00;
      17'd64185: data = 8'h00;
      17'd64186: data = 8'h00;
      17'd64187: data = 8'h01;
      17'd64188: data = 8'h01;
      17'd64189: data = 8'h00;
      17'd64190: data = 8'h01;
      17'd64191: data = 8'h00;
      17'd64192: data = 8'hfe;
      17'd64193: data = 8'hfe;
      17'd64194: data = 8'hfe;
      17'd64195: data = 8'hfe;
      17'd64196: data = 8'hfe;
      17'd64197: data = 8'hfd;
      17'd64198: data = 8'hfe;
      17'd64199: data = 8'hfe;
      17'd64200: data = 8'h01;
      17'd64201: data = 8'h00;
      17'd64202: data = 8'hfe;
      17'd64203: data = 8'h01;
      17'd64204: data = 8'h00;
      17'd64205: data = 8'hfe;
      17'd64206: data = 8'hfe;
      17'd64207: data = 8'h00;
      17'd64208: data = 8'h00;
      17'd64209: data = 8'hfe;
      17'd64210: data = 8'hfe;
      17'd64211: data = 8'hfd;
      17'd64212: data = 8'hfd;
      17'd64213: data = 8'hfe;
      17'd64214: data = 8'hfe;
      17'd64215: data = 8'hfe;
      17'd64216: data = 8'hfe;
      17'd64217: data = 8'hfe;
      17'd64218: data = 8'hfe;
      17'd64219: data = 8'hfe;
      17'd64220: data = 8'hfe;
      17'd64221: data = 8'h00;
      17'd64222: data = 8'hfe;
      17'd64223: data = 8'hfd;
      17'd64224: data = 8'hfd;
      17'd64225: data = 8'hfe;
      17'd64226: data = 8'h00;
      17'd64227: data = 8'hfd;
      17'd64228: data = 8'hfd;
      17'd64229: data = 8'h00;
      17'd64230: data = 8'h01;
      17'd64231: data = 8'h01;
      17'd64232: data = 8'hfe;
      17'd64233: data = 8'hfe;
      17'd64234: data = 8'hfe;
      17'd64235: data = 8'hfd;
      17'd64236: data = 8'hfd;
      17'd64237: data = 8'hfe;
      17'd64238: data = 8'hfd;
      17'd64239: data = 8'hfc;
      17'd64240: data = 8'hfa;
      17'd64241: data = 8'hfc;
      17'd64242: data = 8'hfd;
      17'd64243: data = 8'hfd;
      17'd64244: data = 8'hfe;
      17'd64245: data = 8'hfe;
      17'd64246: data = 8'hfe;
      17'd64247: data = 8'hfd;
      17'd64248: data = 8'hfe;
      17'd64249: data = 8'hfe;
      17'd64250: data = 8'h00;
      17'd64251: data = 8'hfd;
      17'd64252: data = 8'hfa;
      17'd64253: data = 8'hfc;
      17'd64254: data = 8'hfc;
      17'd64255: data = 8'hfa;
      17'd64256: data = 8'hfc;
      17'd64257: data = 8'hfd;
      17'd64258: data = 8'hfd;
      17'd64259: data = 8'hfe;
      17'd64260: data = 8'hfe;
      17'd64261: data = 8'hfe;
      17'd64262: data = 8'hfd;
      17'd64263: data = 8'hfd;
      17'd64264: data = 8'h00;
      17'd64265: data = 8'hfe;
      17'd64266: data = 8'hfe;
      17'd64267: data = 8'hfd;
      17'd64268: data = 8'hfc;
      17'd64269: data = 8'hfc;
      17'd64270: data = 8'hfa;
      17'd64271: data = 8'hfc;
      17'd64272: data = 8'hfd;
      17'd64273: data = 8'hfd;
      17'd64274: data = 8'hfe;
      17'd64275: data = 8'hfe;
      17'd64276: data = 8'hfe;
      17'd64277: data = 8'hfe;
      17'd64278: data = 8'hfe;
      17'd64279: data = 8'hfe;
      17'd64280: data = 8'hfd;
      17'd64281: data = 8'hfe;
      17'd64282: data = 8'hfe;
      17'd64283: data = 8'hfc;
      17'd64284: data = 8'hfd;
      17'd64285: data = 8'hfd;
      17'd64286: data = 8'hfd;
      17'd64287: data = 8'hfd;
      17'd64288: data = 8'hfd;
      17'd64289: data = 8'hfc;
      17'd64290: data = 8'hfe;
      17'd64291: data = 8'hfe;
      17'd64292: data = 8'hfd;
      17'd64293: data = 8'h00;
      17'd64294: data = 8'hfe;
      17'd64295: data = 8'h00;
      17'd64296: data = 8'hfd;
      17'd64297: data = 8'hfc;
      17'd64298: data = 8'hfc;
      17'd64299: data = 8'hfd;
      17'd64300: data = 8'hfd;
      17'd64301: data = 8'hfc;
      17'd64302: data = 8'hfc;
      17'd64303: data = 8'hfd;
      17'd64304: data = 8'hfd;
      17'd64305: data = 8'hfd;
      17'd64306: data = 8'hfd;
      17'd64307: data = 8'hfd;
      17'd64308: data = 8'hfe;
      17'd64309: data = 8'hfe;
      17'd64310: data = 8'hfc;
      17'd64311: data = 8'hfd;
      17'd64312: data = 8'hfd;
      17'd64313: data = 8'hfc;
      17'd64314: data = 8'hfe;
      17'd64315: data = 8'hfe;
      17'd64316: data = 8'hfd;
      17'd64317: data = 8'hfd;
      17'd64318: data = 8'hfd;
      17'd64319: data = 8'hfe;
      17'd64320: data = 8'hfe;
      17'd64321: data = 8'hfe;
      17'd64322: data = 8'hfe;
      17'd64323: data = 8'h00;
      17'd64324: data = 8'h00;
      17'd64325: data = 8'hfe;
      17'd64326: data = 8'hfe;
      17'd64327: data = 8'h01;
      17'd64328: data = 8'h00;
      17'd64329: data = 8'h00;
      17'd64330: data = 8'h00;
      17'd64331: data = 8'hfd;
      17'd64332: data = 8'h00;
      17'd64333: data = 8'h00;
      17'd64334: data = 8'h01;
      17'd64335: data = 8'h01;
      17'd64336: data = 8'h01;
      17'd64337: data = 8'h02;
      17'd64338: data = 8'h01;
      17'd64339: data = 8'h00;
      17'd64340: data = 8'h01;
      17'd64341: data = 8'h02;
      17'd64342: data = 8'h01;
      17'd64343: data = 8'h00;
      17'd64344: data = 8'hfe;
      17'd64345: data = 8'h00;
      17'd64346: data = 8'h00;
      17'd64347: data = 8'h01;
      17'd64348: data = 8'h01;
      17'd64349: data = 8'hfe;
      17'd64350: data = 8'h01;
      17'd64351: data = 8'h01;
      17'd64352: data = 8'h01;
      17'd64353: data = 8'h01;
      17'd64354: data = 8'h01;
      17'd64355: data = 8'h04;
      17'd64356: data = 8'h04;
      17'd64357: data = 8'h02;
      17'd64358: data = 8'h00;
      17'd64359: data = 8'h01;
      17'd64360: data = 8'h00;
      17'd64361: data = 8'h00;
      17'd64362: data = 8'h00;
      17'd64363: data = 8'hfe;
      17'd64364: data = 8'h00;
      17'd64365: data = 8'h00;
      17'd64366: data = 8'h00;
      17'd64367: data = 8'h01;
      17'd64368: data = 8'h02;
      17'd64369: data = 8'h05;
      17'd64370: data = 8'h02;
      17'd64371: data = 8'h02;
      17'd64372: data = 8'h02;
      17'd64373: data = 8'h01;
      17'd64374: data = 8'h00;
      17'd64375: data = 8'h00;
      17'd64376: data = 8'hfe;
      17'd64377: data = 8'hfe;
      17'd64378: data = 8'h01;
      17'd64379: data = 8'h00;
      17'd64380: data = 8'h00;
      17'd64381: data = 8'h01;
      17'd64382: data = 8'h02;
      17'd64383: data = 8'h02;
      17'd64384: data = 8'h04;
      17'd64385: data = 8'h04;
      17'd64386: data = 8'h04;
      17'd64387: data = 8'h04;
      17'd64388: data = 8'h01;
      17'd64389: data = 8'h01;
      17'd64390: data = 8'h01;
      17'd64391: data = 8'h00;
      17'd64392: data = 8'hfe;
      17'd64393: data = 8'hfe;
      17'd64394: data = 8'h00;
      17'd64395: data = 8'h00;
      17'd64396: data = 8'h00;
      17'd64397: data = 8'h01;
      17'd64398: data = 8'h02;
      17'd64399: data = 8'h02;
      17'd64400: data = 8'h02;
      17'd64401: data = 8'h02;
      17'd64402: data = 8'h01;
      17'd64403: data = 8'h01;
      17'd64404: data = 8'h00;
      17'd64405: data = 8'hfe;
      17'd64406: data = 8'hfe;
      17'd64407: data = 8'hfd;
      17'd64408: data = 8'hfc;
      17'd64409: data = 8'hfd;
      17'd64410: data = 8'hfe;
      17'd64411: data = 8'hfe;
      17'd64412: data = 8'h00;
      17'd64413: data = 8'h00;
      17'd64414: data = 8'h01;
      17'd64415: data = 8'h02;
      17'd64416: data = 8'h00;
      17'd64417: data = 8'h04;
      17'd64418: data = 8'h02;
      17'd64419: data = 8'h01;
      17'd64420: data = 8'hfe;
      17'd64421: data = 8'hfe;
      17'd64422: data = 8'h00;
      17'd64423: data = 8'hfc;
      17'd64424: data = 8'hfd;
      17'd64425: data = 8'hfe;
      17'd64426: data = 8'hfe;
      17'd64427: data = 8'h01;
      17'd64428: data = 8'h02;
      17'd64429: data = 8'h01;
      17'd64430: data = 8'h02;
      17'd64431: data = 8'h02;
      17'd64432: data = 8'h01;
      17'd64433: data = 8'h02;
      17'd64434: data = 8'h02;
      17'd64435: data = 8'h01;
      17'd64436: data = 8'hfe;
      17'd64437: data = 8'h00;
      17'd64438: data = 8'h00;
      17'd64439: data = 8'h00;
      17'd64440: data = 8'h02;
      17'd64441: data = 8'h01;
      17'd64442: data = 8'h01;
      17'd64443: data = 8'h02;
      17'd64444: data = 8'h02;
      17'd64445: data = 8'h02;
      17'd64446: data = 8'h04;
      17'd64447: data = 8'h02;
      17'd64448: data = 8'h02;
      17'd64449: data = 8'h00;
      17'd64450: data = 8'h00;
      17'd64451: data = 8'hfe;
      17'd64452: data = 8'hfd;
      17'd64453: data = 8'hfe;
      17'd64454: data = 8'hfe;
      17'd64455: data = 8'h01;
      17'd64456: data = 8'h01;
      17'd64457: data = 8'h01;
      17'd64458: data = 8'h02;
      17'd64459: data = 8'h02;
      17'd64460: data = 8'h02;
      17'd64461: data = 8'h01;
      17'd64462: data = 8'h01;
      17'd64463: data = 8'h01;
      17'd64464: data = 8'hfe;
      17'd64465: data = 8'h00;
      17'd64466: data = 8'h00;
      17'd64467: data = 8'hfe;
      17'd64468: data = 8'hfe;
      17'd64469: data = 8'hfe;
      17'd64470: data = 8'hfe;
      17'd64471: data = 8'h00;
      17'd64472: data = 8'h01;
      17'd64473: data = 8'h00;
      17'd64474: data = 8'h01;
      17'd64475: data = 8'h01;
      17'd64476: data = 8'h00;
      17'd64477: data = 8'hfd;
      17'd64478: data = 8'hfc;
      17'd64479: data = 8'hfd;
      17'd64480: data = 8'hfc;
      17'd64481: data = 8'hfc;
      17'd64482: data = 8'hfd;
      17'd64483: data = 8'hfc;
      17'd64484: data = 8'hfc;
      17'd64485: data = 8'hfd;
      17'd64486: data = 8'hfe;
      17'd64487: data = 8'h00;
      17'd64488: data = 8'h00;
      17'd64489: data = 8'h00;
      17'd64490: data = 8'hfe;
      17'd64491: data = 8'hfe;
      17'd64492: data = 8'hfc;
      17'd64493: data = 8'hfd;
      17'd64494: data = 8'hfc;
      17'd64495: data = 8'hfa;
      17'd64496: data = 8'hfc;
      17'd64497: data = 8'hfd;
      17'd64498: data = 8'hfd;
      17'd64499: data = 8'hfd;
      17'd64500: data = 8'hfd;
      17'd64501: data = 8'hfd;
      17'd64502: data = 8'hfe;
      17'd64503: data = 8'h00;
      17'd64504: data = 8'hfe;
      17'd64505: data = 8'h00;
      17'd64506: data = 8'h00;
      17'd64507: data = 8'hfe;
      17'd64508: data = 8'hfd;
      17'd64509: data = 8'hfd;
      17'd64510: data = 8'hfd;
      17'd64511: data = 8'hfd;
      17'd64512: data = 8'hfd;
      17'd64513: data = 8'hfd;
      17'd64514: data = 8'hfe;
      17'd64515: data = 8'h00;
      17'd64516: data = 8'h00;
      17'd64517: data = 8'h01;
      17'd64518: data = 8'h01;
      17'd64519: data = 8'h00;
      17'd64520: data = 8'h00;
      17'd64521: data = 8'h00;
      17'd64522: data = 8'hfd;
      17'd64523: data = 8'hfd;
      17'd64524: data = 8'hfe;
      17'd64525: data = 8'hfe;
      17'd64526: data = 8'hfe;
      17'd64527: data = 8'hfd;
      17'd64528: data = 8'hfc;
      17'd64529: data = 8'hfd;
      17'd64530: data = 8'hfd;
      17'd64531: data = 8'hfd;
      17'd64532: data = 8'h00;
      17'd64533: data = 8'h01;
      17'd64534: data = 8'h01;
      17'd64535: data = 8'h00;
      17'd64536: data = 8'h01;
      17'd64537: data = 8'h00;
      17'd64538: data = 8'hfe;
      17'd64539: data = 8'hfe;
      17'd64540: data = 8'hfc;
      17'd64541: data = 8'hfd;
      17'd64542: data = 8'hfc;
      17'd64543: data = 8'hfa;
      17'd64544: data = 8'hfc;
      17'd64545: data = 8'hfd;
      17'd64546: data = 8'hfd;
      17'd64547: data = 8'hfe;
      17'd64548: data = 8'h00;
      17'd64549: data = 8'hfd;
      17'd64550: data = 8'hfd;
      17'd64551: data = 8'hfd;
      17'd64552: data = 8'hfc;
      17'd64553: data = 8'hfd;
      17'd64554: data = 8'hfd;
      17'd64555: data = 8'hfc;
      17'd64556: data = 8'hfa;
      17'd64557: data = 8'hfc;
      17'd64558: data = 8'hfc;
      17'd64559: data = 8'hfa;
      17'd64560: data = 8'hfa;
      17'd64561: data = 8'hfa;
      17'd64562: data = 8'hfd;
      17'd64563: data = 8'hfd;
      17'd64564: data = 8'hfc;
      17'd64565: data = 8'hfc;
      17'd64566: data = 8'hfc;
      17'd64567: data = 8'hfd;
      17'd64568: data = 8'hfc;
      17'd64569: data = 8'hfd;
      17'd64570: data = 8'hfc;
      17'd64571: data = 8'hfa;
      17'd64572: data = 8'hfc;
      17'd64573: data = 8'hfc;
      17'd64574: data = 8'hfc;
      17'd64575: data = 8'hfc;
      17'd64576: data = 8'hfe;
      17'd64577: data = 8'hfd;
      17'd64578: data = 8'hfe;
      17'd64579: data = 8'hfe;
      17'd64580: data = 8'hfe;
      17'd64581: data = 8'hfd;
      17'd64582: data = 8'hfd;
      17'd64583: data = 8'hfe;
      17'd64584: data = 8'hfd;
      17'd64585: data = 8'hfd;
      17'd64586: data = 8'hfd;
      17'd64587: data = 8'hfc;
      17'd64588: data = 8'hfc;
      17'd64589: data = 8'hfc;
      17'd64590: data = 8'hfd;
      17'd64591: data = 8'hfe;
      17'd64592: data = 8'hfd;
      17'd64593: data = 8'hfe;
      17'd64594: data = 8'h00;
      17'd64595: data = 8'h00;
      17'd64596: data = 8'h00;
      17'd64597: data = 8'hfe;
      17'd64598: data = 8'hfe;
      17'd64599: data = 8'hfe;
      17'd64600: data = 8'hfe;
      17'd64601: data = 8'h00;
      17'd64602: data = 8'hfe;
      17'd64603: data = 8'hfd;
      17'd64604: data = 8'hfe;
      17'd64605: data = 8'h00;
      17'd64606: data = 8'h00;
      17'd64607: data = 8'h00;
      17'd64608: data = 8'h02;
      17'd64609: data = 8'h02;
      17'd64610: data = 8'h01;
      17'd64611: data = 8'h02;
      17'd64612: data = 8'h04;
      17'd64613: data = 8'h02;
      17'd64614: data = 8'h00;
      17'd64615: data = 8'hfe;
      17'd64616: data = 8'h00;
      17'd64617: data = 8'hfe;
      17'd64618: data = 8'h00;
      17'd64619: data = 8'h01;
      17'd64620: data = 8'h00;
      17'd64621: data = 8'h00;
      17'd64622: data = 8'h02;
      17'd64623: data = 8'h02;
      17'd64624: data = 8'h01;
      17'd64625: data = 8'h02;
      17'd64626: data = 8'h02;
      17'd64627: data = 8'h01;
      17'd64628: data = 8'h01;
      17'd64629: data = 8'h00;
      17'd64630: data = 8'hfe;
      17'd64631: data = 8'h00;
      17'd64632: data = 8'h00;
      17'd64633: data = 8'hfe;
      17'd64634: data = 8'h00;
      17'd64635: data = 8'h02;
      17'd64636: data = 8'h02;
      17'd64637: data = 8'h04;
      17'd64638: data = 8'h04;
      17'd64639: data = 8'h02;
      17'd64640: data = 8'h02;
      17'd64641: data = 8'h02;
      17'd64642: data = 8'h01;
      17'd64643: data = 8'h01;
      17'd64644: data = 8'h01;
      17'd64645: data = 8'hfe;
      17'd64646: data = 8'hfe;
      17'd64647: data = 8'h00;
      17'd64648: data = 8'h00;
      17'd64649: data = 8'h00;
      17'd64650: data = 8'h00;
      17'd64651: data = 8'h00;
      17'd64652: data = 8'h00;
      17'd64653: data = 8'h01;
      17'd64654: data = 8'h02;
      17'd64655: data = 8'h04;
      17'd64656: data = 8'h04;
      17'd64657: data = 8'h01;
      17'd64658: data = 8'h02;
      17'd64659: data = 8'h01;
      17'd64660: data = 8'h00;
      17'd64661: data = 8'hfe;
      17'd64662: data = 8'h00;
      17'd64663: data = 8'hfe;
      17'd64664: data = 8'hfe;
      17'd64665: data = 8'h01;
      17'd64666: data = 8'h01;
      17'd64667: data = 8'h01;
      17'd64668: data = 8'h01;
      17'd64669: data = 8'h02;
      17'd64670: data = 8'h04;
      17'd64671: data = 8'h04;
      17'd64672: data = 8'h02;
      17'd64673: data = 8'h02;
      17'd64674: data = 8'h00;
      17'd64675: data = 8'h01;
      17'd64676: data = 8'h01;
      17'd64677: data = 8'h00;
      17'd64678: data = 8'h00;
      17'd64679: data = 8'h00;
      17'd64680: data = 8'h01;
      17'd64681: data = 8'h00;
      17'd64682: data = 8'h01;
      17'd64683: data = 8'h01;
      17'd64684: data = 8'h04;
      17'd64685: data = 8'h04;
      17'd64686: data = 8'h02;
      17'd64687: data = 8'h05;
      17'd64688: data = 8'h05;
      17'd64689: data = 8'h0a;
      17'd64690: data = 8'h02;
      17'd64691: data = 8'hf2;
      17'd64692: data = 8'hfc;
      17'd64693: data = 8'hfa;
      17'd64694: data = 8'hec;
      17'd64695: data = 8'h01;
      17'd64696: data = 8'h02;
      17'd64697: data = 8'hf9;
      17'd64698: data = 8'h04;
      17'd64699: data = 8'h0a;
      17'd64700: data = 8'h11;
      17'd64701: data = 8'h13;
      17'd64702: data = 8'h0a;
      17'd64703: data = 8'h0a;
      17'd64704: data = 8'h09;
      17'd64705: data = 8'hfe;
      17'd64706: data = 8'hfe;
      17'd64707: data = 8'hf6;
      17'd64708: data = 8'hf4;
      17'd64709: data = 8'hfe;
      17'd64710: data = 8'hfd;
      17'd64711: data = 8'hfa;
      17'd64712: data = 8'h01;
      17'd64713: data = 8'h01;
      17'd64714: data = 8'h01;
      17'd64715: data = 8'h09;
      17'd64716: data = 8'h06;
      17'd64717: data = 8'h09;
      17'd64718: data = 8'h11;
      17'd64719: data = 8'h0d;
      17'd64720: data = 8'h0e;
      17'd64721: data = 8'hfd;
      17'd64722: data = 8'hef;
      17'd64723: data = 8'hef;
      17'd64724: data = 8'he7;
      17'd64725: data = 8'he9;
      17'd64726: data = 8'heb;
      17'd64727: data = 8'hf4;
      17'd64728: data = 8'hfe;
      17'd64729: data = 8'h0d;
      17'd64730: data = 8'h12;
      17'd64731: data = 8'h0d;
      17'd64732: data = 8'h0a;
      17'd64733: data = 8'h02;
      17'd64734: data = 8'hfc;
      17'd64735: data = 8'hef;
      17'd64736: data = 8'hec;
      17'd64737: data = 8'he5;
      17'd64738: data = 8'he5;
      17'd64739: data = 8'hef;
      17'd64740: data = 8'hf2;
      17'd64741: data = 8'hfc;
      17'd64742: data = 8'hfe;
      17'd64743: data = 8'h09;
      17'd64744: data = 8'h0c;
      17'd64745: data = 8'h0c;
      17'd64746: data = 8'h0c;
      17'd64747: data = 8'h09;
      17'd64748: data = 8'h05;
      17'd64749: data = 8'h01;
      17'd64750: data = 8'hfd;
      17'd64751: data = 8'hf4;
      17'd64752: data = 8'hf1;
      17'd64753: data = 8'hf4;
      17'd64754: data = 8'hf5;
      17'd64755: data = 8'hfa;
      17'd64756: data = 8'h01;
      17'd64757: data = 8'h04;
      17'd64758: data = 8'h09;
      17'd64759: data = 8'h0d;
      17'd64760: data = 8'h0e;
      17'd64761: data = 8'h0e;
      17'd64762: data = 8'h0c;
      17'd64763: data = 8'h05;
      17'd64764: data = 8'hfe;
      17'd64765: data = 8'hf9;
      17'd64766: data = 8'hf9;
      17'd64767: data = 8'hfa;
      17'd64768: data = 8'hfc;
      17'd64769: data = 8'hfe;
      17'd64770: data = 8'h02;
      17'd64771: data = 8'h06;
      17'd64772: data = 8'h09;
      17'd64773: data = 8'h09;
      17'd64774: data = 8'h05;
      17'd64775: data = 8'h05;
      17'd64776: data = 8'h01;
      17'd64777: data = 8'h00;
      17'd64778: data = 8'h00;
      17'd64779: data = 8'hfc;
      17'd64780: data = 8'hfa;
      17'd64781: data = 8'hfa;
      17'd64782: data = 8'hfc;
      17'd64783: data = 8'h00;
      17'd64784: data = 8'h01;
      17'd64785: data = 8'h01;
      17'd64786: data = 8'h04;
      17'd64787: data = 8'h00;
      17'd64788: data = 8'h00;
      17'd64789: data = 8'hfc;
      17'd64790: data = 8'hfa;
      17'd64791: data = 8'hfa;
      17'd64792: data = 8'hf5;
      17'd64793: data = 8'hf9;
      17'd64794: data = 8'hfa;
      17'd64795: data = 8'hf9;
      17'd64796: data = 8'hfd;
      17'd64797: data = 8'h00;
      17'd64798: data = 8'h00;
      17'd64799: data = 8'h00;
      17'd64800: data = 8'hfe;
      17'd64801: data = 8'hfa;
      17'd64802: data = 8'hf9;
      17'd64803: data = 8'hf4;
      17'd64804: data = 8'hf2;
      17'd64805: data = 8'hf5;
      17'd64806: data = 8'hf6;
      17'd64807: data = 8'hf9;
      17'd64808: data = 8'hf9;
      17'd64809: data = 8'hfd;
      17'd64810: data = 8'hfe;
      17'd64811: data = 8'hfe;
      17'd64812: data = 8'hfd;
      17'd64813: data = 8'hfd;
      17'd64814: data = 8'hfc;
      17'd64815: data = 8'hfc;
      17'd64816: data = 8'hfa;
      17'd64817: data = 8'hf9;
      17'd64818: data = 8'hf6;
      17'd64819: data = 8'hf5;
      17'd64820: data = 8'hf9;
      17'd64821: data = 8'hf9;
      17'd64822: data = 8'hfa;
      17'd64823: data = 8'hfe;
      17'd64824: data = 8'hfd;
      17'd64825: data = 8'hfe;
      17'd64826: data = 8'h00;
      17'd64827: data = 8'h00;
      17'd64828: data = 8'h00;
      17'd64829: data = 8'hfe;
      17'd64830: data = 8'hfd;
      17'd64831: data = 8'hfd;
      17'd64832: data = 8'hf9;
      17'd64833: data = 8'hf9;
      17'd64834: data = 8'hf9;
      17'd64835: data = 8'hf9;
      17'd64836: data = 8'hf9;
      17'd64837: data = 8'hfd;
      17'd64838: data = 8'h00;
      17'd64839: data = 8'h00;
      17'd64840: data = 8'h00;
      17'd64841: data = 8'h01;
      17'd64842: data = 8'h02;
      17'd64843: data = 8'h04;
      17'd64844: data = 8'h05;
      17'd64845: data = 8'hfe;
      17'd64846: data = 8'hfd;
      17'd64847: data = 8'hfa;
      17'd64848: data = 8'hf5;
      17'd64849: data = 8'hf4;
      17'd64850: data = 8'hf6;
      17'd64851: data = 8'hf5;
      17'd64852: data = 8'h02;
      17'd64853: data = 8'h06;
      17'd64854: data = 8'h05;
      17'd64855: data = 8'h09;
      17'd64856: data = 8'h01;
      17'd64857: data = 8'h00;
      17'd64858: data = 8'h01;
      17'd64859: data = 8'hfa;
      17'd64860: data = 8'hf9;
      17'd64861: data = 8'hf5;
      17'd64862: data = 8'hf5;
      17'd64863: data = 8'hfd;
      17'd64864: data = 8'h00;
      17'd64865: data = 8'h04;
      17'd64866: data = 8'h04;
      17'd64867: data = 8'h05;
      17'd64868: data = 8'h02;
      17'd64869: data = 8'hfc;
      17'd64870: data = 8'hfc;
      17'd64871: data = 8'hfa;
      17'd64872: data = 8'hfa;
      17'd64873: data = 8'h00;
      17'd64874: data = 8'h02;
      17'd64875: data = 8'h06;
      17'd64876: data = 8'h06;
      17'd64877: data = 8'h02;
      17'd64878: data = 8'h00;
      17'd64879: data = 8'hfa;
      17'd64880: data = 8'hfd;
      17'd64881: data = 8'hfd;
      17'd64882: data = 8'h00;
      17'd64883: data = 8'h04;
      17'd64884: data = 8'h05;
      17'd64885: data = 8'h05;
      17'd64886: data = 8'h00;
      17'd64887: data = 8'h00;
      17'd64888: data = 8'h02;
      17'd64889: data = 8'h01;
      17'd64890: data = 8'hf9;
      17'd64891: data = 8'hfc;
      17'd64892: data = 8'h01;
      17'd64893: data = 8'hfe;
      17'd64894: data = 8'h04;
      17'd64895: data = 8'h06;
      17'd64896: data = 8'h09;
      17'd64897: data = 8'h06;
      17'd64898: data = 8'h02;
      17'd64899: data = 8'h02;
      17'd64900: data = 8'hfe;
      17'd64901: data = 8'hfe;
      17'd64902: data = 8'hfe;
      17'd64903: data = 8'hfc;
      17'd64904: data = 8'h00;
      17'd64905: data = 8'h05;
      17'd64906: data = 8'h06;
      17'd64907: data = 8'h0a;
      17'd64908: data = 8'h0e;
      17'd64909: data = 8'h01;
      17'd64910: data = 8'h05;
      17'd64911: data = 8'h06;
      17'd64912: data = 8'h00;
      17'd64913: data = 8'h00;
      17'd64914: data = 8'h00;
      17'd64915: data = 8'hfe;
      17'd64916: data = 8'h00;
      17'd64917: data = 8'h00;
      17'd64918: data = 8'h01;
      17'd64919: data = 8'h04;
      17'd64920: data = 8'h04;
      17'd64921: data = 8'h0c;
      17'd64922: data = 8'h05;
      17'd64923: data = 8'h01;
      17'd64924: data = 8'hfa;
      17'd64925: data = 8'hf6;
      17'd64926: data = 8'hfc;
      17'd64927: data = 8'hfd;
      17'd64928: data = 8'h01;
      17'd64929: data = 8'h06;
      17'd64930: data = 8'h0c;
      17'd64931: data = 8'h0c;
      17'd64932: data = 8'h0a;
      17'd64933: data = 8'hfe;
      17'd64934: data = 8'hfa;
      17'd64935: data = 8'hf4;
      17'd64936: data = 8'he7;
      17'd64937: data = 8'hed;
      17'd64938: data = 8'hf5;
      17'd64939: data = 8'h02;
      17'd64940: data = 8'h11;
      17'd64941: data = 8'h1e;
      17'd64942: data = 8'h1a;
      17'd64943: data = 8'h06;
      17'd64944: data = 8'hfa;
      17'd64945: data = 8'he9;
      17'd64946: data = 8'he3;
      17'd64947: data = 8'he7;
      17'd64948: data = 8'hf6;
      17'd64949: data = 8'h02;
      17'd64950: data = 8'h05;
      17'd64951: data = 8'h15;
      17'd64952: data = 8'h1a;
      17'd64953: data = 8'h0a;
      17'd64954: data = 8'h00;
      17'd64955: data = 8'hf2;
      17'd64956: data = 8'hf2;
      17'd64957: data = 8'hf1;
      17'd64958: data = 8'hf2;
      17'd64959: data = 8'h00;
      17'd64960: data = 8'h05;
      17'd64961: data = 8'h0e;
      17'd64962: data = 8'h11;
      17'd64963: data = 8'h12;
      17'd64964: data = 8'h0a;
      17'd64965: data = 8'hf5;
      17'd64966: data = 8'hef;
      17'd64967: data = 8'hec;
      17'd64968: data = 8'hfa;
      17'd64969: data = 8'h00;
      17'd64970: data = 8'h04;
      17'd64971: data = 8'h0c;
      17'd64972: data = 8'h0a;
      17'd64973: data = 8'h09;
      17'd64974: data = 8'h00;
      17'd64975: data = 8'hfe;
      17'd64976: data = 8'hfc;
      17'd64977: data = 8'hfa;
      17'd64978: data = 8'hfe;
      17'd64979: data = 8'h02;
      17'd64980: data = 8'h05;
      17'd64981: data = 8'h0a;
      17'd64982: data = 8'h06;
      17'd64983: data = 8'h11;
      17'd64984: data = 8'h02;
      17'd64985: data = 8'hf2;
      17'd64986: data = 8'hfa;
      17'd64987: data = 8'hed;
      17'd64988: data = 8'hef;
      17'd64989: data = 8'hfd;
      17'd64990: data = 8'h05;
      17'd64991: data = 8'h13;
      17'd64992: data = 8'h12;
      17'd64993: data = 8'h0e;
      17'd64994: data = 8'h04;
      17'd64995: data = 8'hf9;
      17'd64996: data = 8'hf5;
      17'd64997: data = 8'hed;
      17'd64998: data = 8'hec;
      17'd64999: data = 8'hef;
      17'd65000: data = 8'hf6;
      17'd65001: data = 8'h01;
      17'd65002: data = 8'h15;
      17'd65003: data = 8'h0a;
      17'd65004: data = 8'h02;
      17'd65005: data = 8'hfe;
      17'd65006: data = 8'hf4;
      17'd65007: data = 8'h00;
      17'd65008: data = 8'hef;
      17'd65009: data = 8'hed;
      17'd65010: data = 8'hfc;
      17'd65011: data = 8'h01;
      17'd65012: data = 8'h0c;
      17'd65013: data = 8'h06;
      17'd65014: data = 8'h04;
      17'd65015: data = 8'h04;
      17'd65016: data = 8'hf5;
      17'd65017: data = 8'hf1;
      17'd65018: data = 8'hf4;
      17'd65019: data = 8'hf4;
      17'd65020: data = 8'hf6;
      17'd65021: data = 8'h05;
      17'd65022: data = 8'h01;
      17'd65023: data = 8'h05;
      17'd65024: data = 8'h0e;
      17'd65025: data = 8'hfc;
      17'd65026: data = 8'hfe;
      17'd65027: data = 8'h00;
      17'd65028: data = 8'hf9;
      17'd65029: data = 8'hf4;
      17'd65030: data = 8'hf2;
      17'd65031: data = 8'hfe;
      17'd65032: data = 8'hfd;
      17'd65033: data = 8'h02;
      17'd65034: data = 8'h0d;
      17'd65035: data = 8'h0c;
      17'd65036: data = 8'h04;
      17'd65037: data = 8'hfd;
      17'd65038: data = 8'hfc;
      17'd65039: data = 8'hf1;
      17'd65040: data = 8'hf4;
      17'd65041: data = 8'hfd;
      17'd65042: data = 8'hf6;
      17'd65043: data = 8'hfe;
      17'd65044: data = 8'h0a;
      17'd65045: data = 8'h0c;
      17'd65046: data = 8'h0a;
      17'd65047: data = 8'hfc;
      17'd65048: data = 8'h00;
      17'd65049: data = 8'hfd;
      17'd65050: data = 8'hf4;
      17'd65051: data = 8'hfa;
      17'd65052: data = 8'hfa;
      17'd65053: data = 8'hfe;
      17'd65054: data = 8'h04;
      17'd65055: data = 8'h02;
      17'd65056: data = 8'h0c;
      17'd65057: data = 8'h06;
      17'd65058: data = 8'hfa;
      17'd65059: data = 8'h01;
      17'd65060: data = 8'hfd;
      17'd65061: data = 8'hf5;
      17'd65062: data = 8'h02;
      17'd65063: data = 8'h06;
      17'd65064: data = 8'hf9;
      17'd65065: data = 8'hfc;
      17'd65066: data = 8'h01;
      17'd65067: data = 8'h04;
      17'd65068: data = 8'h04;
      17'd65069: data = 8'h09;
      17'd65070: data = 8'h05;
      17'd65071: data = 8'hf5;
      17'd65072: data = 8'hfd;
      17'd65073: data = 8'h02;
      17'd65074: data = 8'h01;
      17'd65075: data = 8'h00;
      17'd65076: data = 8'h09;
      17'd65077: data = 8'h04;
      17'd65078: data = 8'hf6;
      17'd65079: data = 8'hfe;
      17'd65080: data = 8'h02;
      17'd65081: data = 8'hf9;
      17'd65082: data = 8'hfa;
      17'd65083: data = 8'h05;
      17'd65084: data = 8'h05;
      17'd65085: data = 8'h06;
      17'd65086: data = 8'h06;
      17'd65087: data = 8'h09;
      17'd65088: data = 8'hfe;
      17'd65089: data = 8'hf5;
      17'd65090: data = 8'hfa;
      17'd65091: data = 8'hfc;
      17'd65092: data = 8'hf9;
      17'd65093: data = 8'h04;
      17'd65094: data = 8'h04;
      17'd65095: data = 8'h02;
      17'd65096: data = 8'h09;
      17'd65097: data = 8'h04;
      17'd65098: data = 8'h04;
      17'd65099: data = 8'hfe;
      17'd65100: data = 8'hf6;
      17'd65101: data = 8'hf9;
      17'd65102: data = 8'hfa;
      17'd65103: data = 8'hfc;
      17'd65104: data = 8'h00;
      17'd65105: data = 8'h02;
      17'd65106: data = 8'h02;
      17'd65107: data = 8'h01;
      17'd65108: data = 8'h00;
      17'd65109: data = 8'hf9;
      17'd65110: data = 8'hf5;
      17'd65111: data = 8'hfc;
      17'd65112: data = 8'hfd;
      17'd65113: data = 8'hfa;
      17'd65114: data = 8'hfd;
      17'd65115: data = 8'h00;
      17'd65116: data = 8'hfc;
      17'd65117: data = 8'hfd;
      17'd65118: data = 8'hfc;
      17'd65119: data = 8'hf9;
      17'd65120: data = 8'hf9;
      17'd65121: data = 8'hfa;
      17'd65122: data = 8'hfa;
      17'd65123: data = 8'hfe;
      17'd65124: data = 8'h01;
      17'd65125: data = 8'hfe;
      17'd65126: data = 8'hfa;
      17'd65127: data = 8'hfd;
      17'd65128: data = 8'hfa;
      17'd65129: data = 8'hf1;
      17'd65130: data = 8'hf2;
      17'd65131: data = 8'hfe;
      17'd65132: data = 8'hfd;
      17'd65133: data = 8'h01;
      17'd65134: data = 8'h05;
      17'd65135: data = 8'h02;
      17'd65136: data = 8'h02;
      17'd65137: data = 8'hf9;
      17'd65138: data = 8'hf6;
      17'd65139: data = 8'hf2;
      17'd65140: data = 8'hf4;
      17'd65141: data = 8'hfc;
      17'd65142: data = 8'hfe;
      17'd65143: data = 8'h02;
      17'd65144: data = 8'h0a;
      17'd65145: data = 8'h0a;
      17'd65146: data = 8'h06;
      17'd65147: data = 8'h09;
      17'd65148: data = 8'hfd;
      17'd65149: data = 8'hf4;
      17'd65150: data = 8'hf5;
      17'd65151: data = 8'hf4;
      17'd65152: data = 8'hfc;
      17'd65153: data = 8'h05;
      17'd65154: data = 8'h0e;
      17'd65155: data = 8'h12;
      17'd65156: data = 8'h0a;
      17'd65157: data = 8'h04;
      17'd65158: data = 8'h02;
      17'd65159: data = 8'h02;
      17'd65160: data = 8'h01;
      17'd65161: data = 8'h00;
      17'd65162: data = 8'hfd;
      17'd65163: data = 8'h01;
      17'd65164: data = 8'h04;
      17'd65165: data = 8'h05;
      17'd65166: data = 8'h0a;
      17'd65167: data = 8'h0e;
      17'd65168: data = 8'h0c;
      17'd65169: data = 8'h04;
      17'd65170: data = 8'h06;
      17'd65171: data = 8'h01;
      17'd65172: data = 8'h01;
      17'd65173: data = 8'hfe;
      17'd65174: data = 8'h01;
      17'd65175: data = 8'h09;
      17'd65176: data = 8'h05;
      17'd65177: data = 8'h09;
      17'd65178: data = 8'h06;
      17'd65179: data = 8'h02;
      17'd65180: data = 8'h04;
      17'd65181: data = 8'h01;
      17'd65182: data = 8'hfc;
      17'd65183: data = 8'h05;
      17'd65184: data = 8'h04;
      17'd65185: data = 8'h06;
      17'd65186: data = 8'h06;
      17'd65187: data = 8'hfa;
      17'd65188: data = 8'h00;
      17'd65189: data = 8'h00;
      17'd65190: data = 8'h00;
      17'd65191: data = 8'h04;
      17'd65192: data = 8'h00;
      17'd65193: data = 8'hfc;
      17'd65194: data = 8'hfd;
      17'd65195: data = 8'hfd;
      17'd65196: data = 8'hfa;
      17'd65197: data = 8'hfd;
      17'd65198: data = 8'h02;
      17'd65199: data = 8'h05;
      17'd65200: data = 8'hfc;
      17'd65201: data = 8'hfd;
      17'd65202: data = 8'hfc;
      17'd65203: data = 8'hef;
      17'd65204: data = 8'hf1;
      17'd65205: data = 8'hfe;
      17'd65206: data = 8'hf6;
      17'd65207: data = 8'hf5;
      17'd65208: data = 8'h04;
      17'd65209: data = 8'hfd;
      17'd65210: data = 8'hf4;
      17'd65211: data = 8'hef;
      17'd65212: data = 8'hf4;
      17'd65213: data = 8'hfc;
      17'd65214: data = 8'hf9;
      17'd65215: data = 8'hf5;
      17'd65216: data = 8'h01;
      17'd65217: data = 8'hf9;
      17'd65218: data = 8'hfe;
      17'd65219: data = 8'h01;
      17'd65220: data = 8'hef;
      17'd65221: data = 8'hec;
      17'd65222: data = 8'hf6;
      17'd65223: data = 8'hf5;
      17'd65224: data = 8'hf1;
      17'd65225: data = 8'h00;
      17'd65226: data = 8'h00;
      17'd65227: data = 8'h00;
      17'd65228: data = 8'h04;
      17'd65229: data = 8'h00;
      17'd65230: data = 8'hfa;
      17'd65231: data = 8'heb;
      17'd65232: data = 8'hf2;
      17'd65233: data = 8'h01;
      17'd65234: data = 8'hf2;
      17'd65235: data = 8'h09;
      17'd65236: data = 8'h12;
      17'd65237: data = 8'h0c;
      17'd65238: data = 8'h1a;
      17'd65239: data = 8'hfc;
      17'd65240: data = 8'hf4;
      17'd65241: data = 8'hf1;
      17'd65242: data = 8'hf1;
      17'd65243: data = 8'h00;
      17'd65244: data = 8'hfe;
      17'd65245: data = 8'h09;
      17'd65246: data = 8'h0c;
      17'd65247: data = 8'h11;
      17'd65248: data = 8'h0a;
      17'd65249: data = 8'h06;
      17'd65250: data = 8'h05;
      17'd65251: data = 8'hfa;
      17'd65252: data = 8'h06;
      17'd65253: data = 8'h09;
      17'd65254: data = 8'h00;
      17'd65255: data = 8'hfc;
      17'd65256: data = 8'h00;
      17'd65257: data = 8'h0a;
      17'd65258: data = 8'h09;
      17'd65259: data = 8'h02;
      17'd65260: data = 8'h02;
      17'd65261: data = 8'hfd;
      17'd65262: data = 8'hfc;
      17'd65263: data = 8'h00;
      17'd65264: data = 8'hfd;
      17'd65265: data = 8'h04;
      17'd65266: data = 8'h12;
      17'd65267: data = 8'h0e;
      17'd65268: data = 8'h02;
      17'd65269: data = 8'hf5;
      17'd65270: data = 8'hf1;
      17'd65271: data = 8'h00;
      17'd65272: data = 8'h02;
      17'd65273: data = 8'h02;
      17'd65274: data = 8'h0e;
      17'd65275: data = 8'h0c;
      17'd65276: data = 8'h04;
      17'd65277: data = 8'h00;
      17'd65278: data = 8'hf5;
      17'd65279: data = 8'hf9;
      17'd65280: data = 8'hf4;
      17'd65281: data = 8'hf4;
      17'd65282: data = 8'h02;
      17'd65283: data = 8'h05;
      17'd65284: data = 8'h09;
      17'd65285: data = 8'h0a;
      17'd65286: data = 8'h06;
      17'd65287: data = 8'h01;
      17'd65288: data = 8'h00;
      17'd65289: data = 8'hfa;
      17'd65290: data = 8'hf6;
      17'd65291: data = 8'hfc;
      17'd65292: data = 8'hf6;
      17'd65293: data = 8'hfa;
      17'd65294: data = 8'h05;
      17'd65295: data = 8'h09;
      17'd65296: data = 8'h09;
      17'd65297: data = 8'h02;
      17'd65298: data = 8'hf2;
      17'd65299: data = 8'hf1;
      17'd65300: data = 8'hf6;
      17'd65301: data = 8'h00;
      17'd65302: data = 8'h05;
      17'd65303: data = 8'h04;
      17'd65304: data = 8'h05;
      17'd65305: data = 8'h04;
      17'd65306: data = 8'hfa;
      17'd65307: data = 8'hfc;
      17'd65308: data = 8'hfc;
      17'd65309: data = 8'hf6;
      17'd65310: data = 8'h01;
      17'd65311: data = 8'h04;
      17'd65312: data = 8'h02;
      17'd65313: data = 8'h09;
      17'd65314: data = 8'h09;
      17'd65315: data = 8'h05;
      17'd65316: data = 8'h02;
      17'd65317: data = 8'hfc;
      17'd65318: data = 8'hfe;
      17'd65319: data = 8'hfd;
      17'd65320: data = 8'hfd;
      17'd65321: data = 8'h04;
      17'd65322: data = 8'h04;
      17'd65323: data = 8'h05;
      17'd65324: data = 8'h0c;
      17'd65325: data = 8'h0c;
      17'd65326: data = 8'h02;
      17'd65327: data = 8'hfe;
      17'd65328: data = 8'hfc;
      17'd65329: data = 8'hfe;
      17'd65330: data = 8'h05;
      17'd65331: data = 8'h0d;
      17'd65332: data = 8'h0d;
      17'd65333: data = 8'h06;
      17'd65334: data = 8'h01;
      17'd65335: data = 8'hfd;
      17'd65336: data = 8'hf9;
      17'd65337: data = 8'hfd;
      17'd65338: data = 8'h02;
      17'd65339: data = 8'h01;
      17'd65340: data = 8'h02;
      17'd65341: data = 8'h06;
      17'd65342: data = 8'h04;
      17'd65343: data = 8'h01;
      17'd65344: data = 8'h02;
      17'd65345: data = 8'hfd;
      17'd65346: data = 8'hf9;
      17'd65347: data = 8'hfa;
      17'd65348: data = 8'hf9;
      17'd65349: data = 8'hfd;
      17'd65350: data = 8'hfd;
      17'd65351: data = 8'hfa;
      17'd65352: data = 8'hfa;
      17'd65353: data = 8'hf9;
      17'd65354: data = 8'hf9;
      17'd65355: data = 8'hf5;
      17'd65356: data = 8'hf5;
      17'd65357: data = 8'hf4;
      17'd65358: data = 8'hf5;
      17'd65359: data = 8'hf9;
      17'd65360: data = 8'hfa;
      17'd65361: data = 8'hf9;
      17'd65362: data = 8'hf6;
      17'd65363: data = 8'hf5;
      17'd65364: data = 8'hf2;
      17'd65365: data = 8'hf4;
      17'd65366: data = 8'hf5;
      17'd65367: data = 8'hf5;
      17'd65368: data = 8'hfa;
      17'd65369: data = 8'hf9;
      17'd65370: data = 8'hf9;
      17'd65371: data = 8'hf6;
      17'd65372: data = 8'hfa;
      17'd65373: data = 8'hfc;
      17'd65374: data = 8'hfe;
      17'd65375: data = 8'hfe;
      17'd65376: data = 8'hfc;
      17'd65377: data = 8'hfd;
      17'd65378: data = 8'hfd;
      17'd65379: data = 8'h00;
      17'd65380: data = 8'h00;
      17'd65381: data = 8'h01;
      17'd65382: data = 8'h01;
      17'd65383: data = 8'hfe;
      17'd65384: data = 8'hfd;
      17'd65385: data = 8'h01;
      17'd65386: data = 8'h02;
      17'd65387: data = 8'h05;
      17'd65388: data = 8'h06;
      17'd65389: data = 8'h09;
      17'd65390: data = 8'h09;
      17'd65391: data = 8'h05;
      17'd65392: data = 8'h04;
      17'd65393: data = 8'h01;
      17'd65394: data = 8'h02;
      17'd65395: data = 8'h02;
      17'd65396: data = 8'h04;
      17'd65397: data = 8'h05;
      17'd65398: data = 8'h06;
      17'd65399: data = 8'h09;
      17'd65400: data = 8'h09;
      17'd65401: data = 8'h0a;
      17'd65402: data = 8'h06;
      17'd65403: data = 8'h05;
      17'd65404: data = 8'h02;
      17'd65405: data = 8'hfe;
      17'd65406: data = 8'h01;
      17'd65407: data = 8'h04;
      17'd65408: data = 8'h06;
      17'd65409: data = 8'h0a;
      17'd65410: data = 8'h0a;
      17'd65411: data = 8'h04;
      17'd65412: data = 8'h00;
      17'd65413: data = 8'h01;
      17'd65414: data = 8'hfd;
      17'd65415: data = 8'hfe;
      17'd65416: data = 8'h06;
      17'd65417: data = 8'h06;
      17'd65418: data = 8'h06;
      17'd65419: data = 8'h0a;
      17'd65420: data = 8'h05;
      17'd65421: data = 8'h01;
      17'd65422: data = 8'hfe;
      17'd65423: data = 8'hf9;
      17'd65424: data = 8'hf5;
      17'd65425: data = 8'hf6;
      17'd65426: data = 8'hfc;
      17'd65427: data = 8'hfa;
      17'd65428: data = 8'hfc;
      17'd65429: data = 8'h01;
      17'd65430: data = 8'h00;
      17'd65431: data = 8'hfd;
      17'd65432: data = 8'hfc;
      17'd65433: data = 8'hf6;
      17'd65434: data = 8'hf4;
      17'd65435: data = 8'hf6;
      17'd65436: data = 8'hf6;
      17'd65437: data = 8'hfa;
      17'd65438: data = 8'hfc;
      17'd65439: data = 8'hf9;
      17'd65440: data = 8'hf9;
      17'd65441: data = 8'hf9;
      17'd65442: data = 8'hf4;
      17'd65443: data = 8'hf5;
      17'd65444: data = 8'hf6;
      17'd65445: data = 8'hf4;
      17'd65446: data = 8'hf4;
      17'd65447: data = 8'hf9;
      17'd65448: data = 8'hfc;
      17'd65449: data = 8'hf4;
      17'd65450: data = 8'hf4;
      17'd65451: data = 8'hf4;
      17'd65452: data = 8'hef;
      17'd65453: data = 8'hf5;
      17'd65454: data = 8'hf6;
      17'd65455: data = 8'hf9;
      17'd65456: data = 8'hf9;
      17'd65457: data = 8'hf9;
      17'd65458: data = 8'hfa;
      17'd65459: data = 8'hf1;
      17'd65460: data = 8'hf5;
      17'd65461: data = 8'hf5;
      17'd65462: data = 8'hed;
      17'd65463: data = 8'hf5;
      17'd65464: data = 8'hfa;
      17'd65465: data = 8'h00;
      17'd65466: data = 8'hfe;
      17'd65467: data = 8'hfe;
      17'd65468: data = 8'hf6;
      17'd65469: data = 8'hf1;
      17'd65470: data = 8'hf5;
      17'd65471: data = 8'hf4;
      17'd65472: data = 8'hfc;
      17'd65473: data = 8'h01;
      17'd65474: data = 8'h00;
      17'd65475: data = 8'h00;
      17'd65476: data = 8'h00;
      17'd65477: data = 8'h00;
      17'd65478: data = 8'h06;
      17'd65479: data = 8'h05;
      17'd65480: data = 8'hfe;
      17'd65481: data = 8'hf6;
      17'd65482: data = 8'hfe;
      17'd65483: data = 8'h06;
      17'd65484: data = 8'h05;
      17'd65485: data = 8'h0e;
      17'd65486: data = 8'h06;
      17'd65487: data = 8'h01;
      17'd65488: data = 8'h05;
      17'd65489: data = 8'h05;
      17'd65490: data = 8'h0c;
      17'd65491: data = 8'h09;
      17'd65492: data = 8'h04;
      17'd65493: data = 8'h0c;
      17'd65494: data = 8'h04;
      17'd65495: data = 8'h0d;
      17'd65496: data = 8'h15;
      17'd65497: data = 8'h09;
      17'd65498: data = 8'h0c;
      17'd65499: data = 8'h0d;
      17'd65500: data = 8'h0a;
      17'd65501: data = 8'h0e;
      17'd65502: data = 8'h0d;
      17'd65503: data = 8'h02;
      17'd65504: data = 8'h01;
      17'd65505: data = 8'h04;
      17'd65506: data = 8'h0c;
      17'd65507: data = 8'h0a;
      17'd65508: data = 8'h0e;
      17'd65509: data = 8'h1b;
      17'd65510: data = 8'h11;
      17'd65511: data = 8'h05;
      17'd65512: data = 8'h01;
      17'd65513: data = 8'h02;
      17'd65514: data = 8'h00;
      17'd65515: data = 8'h01;
      17'd65516: data = 8'h05;
      17'd65517: data = 8'h0c;
      17'd65518: data = 8'h12;
      17'd65519: data = 8'h09;
      17'd65520: data = 8'h0a;
      17'd65521: data = 8'h02;
      17'd65522: data = 8'hf4;
      17'd65523: data = 8'h00;
      17'd65524: data = 8'hfe;
      17'd65525: data = 8'hfa;
      17'd65526: data = 8'h0d;
      17'd65527: data = 8'h0c;
      17'd65528: data = 8'hfc;
      17'd65529: data = 8'h04;
      17'd65530: data = 8'h0e;
      17'd65531: data = 8'hfc;
      17'd65532: data = 8'hef;
      17'd65533: data = 8'hfa;
      17'd65534: data = 8'hf2;
      17'd65535: data = 8'hf4;
      17'd65536: data = 8'h05;
      17'd65537: data = 8'h09;
      17'd65538: data = 8'h09;
      17'd65539: data = 8'h06;
      17'd65540: data = 8'h04;
      17'd65541: data = 8'hf9;
      17'd65542: data = 8'he9;
      17'd65543: data = 8'hf1;
      17'd65544: data = 8'hfd;
      17'd65545: data = 8'h00;
      17'd65546: data = 8'h09;
      17'd65547: data = 8'h0e;
      17'd65548: data = 8'h04;
      17'd65549: data = 8'h04;
      17'd65550: data = 8'hfd;
      17'd65551: data = 8'hf4;
      17'd65552: data = 8'hf1;
      17'd65553: data = 8'hf5;
      17'd65554: data = 8'hfe;
      17'd65555: data = 8'hfd;
      17'd65556: data = 8'h05;
      17'd65557: data = 8'h06;
      17'd65558: data = 8'hfd;
      17'd65559: data = 8'h00;
      17'd65560: data = 8'h04;
      17'd65561: data = 8'hfe;
      17'd65562: data = 8'hf9;
      17'd65563: data = 8'hf5;
      17'd65564: data = 8'hf5;
      17'd65565: data = 8'hf4;
      17'd65566: data = 8'h01;
      17'd65567: data = 8'h09;
      17'd65568: data = 8'h02;
      17'd65569: data = 8'h09;
      17'd65570: data = 8'h00;
      17'd65571: data = 8'hf5;
      17'd65572: data = 8'hfa;
      17'd65573: data = 8'h00;
      17'd65574: data = 8'h06;
      17'd65575: data = 8'h0a;
      17'd65576: data = 8'h04;
      17'd65577: data = 8'hfa;
      17'd65578: data = 8'hf6;
      17'd65579: data = 8'hfa;
      17'd65580: data = 8'hfa;
      17'd65581: data = 8'h00;
      17'd65582: data = 8'h0a;
      17'd65583: data = 8'h0c;
      17'd65584: data = 8'h04;
      17'd65585: data = 8'h02;
      17'd65586: data = 8'hfd;
      17'd65587: data = 8'hf9;
      17'd65588: data = 8'h01;
      17'd65589: data = 8'h06;
      17'd65590: data = 8'h02;
      17'd65591: data = 8'h00;
      17'd65592: data = 8'h01;
      17'd65593: data = 8'hf4;
      17'd65594: data = 8'hf6;
      17'd65595: data = 8'h04;
      17'd65596: data = 8'h04;
      17'd65597: data = 8'h05;
      17'd65598: data = 8'h04;
      17'd65599: data = 8'hf9;
      17'd65600: data = 8'hf2;
      17'd65601: data = 8'hf4;
      17'd65602: data = 8'hf6;
      17'd65603: data = 8'hfd;
      17'd65604: data = 8'h01;
      17'd65605: data = 8'h00;
      17'd65606: data = 8'hf2;
      17'd65607: data = 8'hef;
      17'd65608: data = 8'hf2;
      17'd65609: data = 8'hf4;
      17'd65610: data = 8'hf9;
      17'd65611: data = 8'hfc;
      17'd65612: data = 8'hf6;
      17'd65613: data = 8'hed;
      17'd65614: data = 8'hec;
      17'd65615: data = 8'he9;
      17'd65616: data = 8'hed;
      17'd65617: data = 8'hf6;
      17'd65618: data = 8'hfc;
      17'd65619: data = 8'hfc;
      17'd65620: data = 8'hf4;
      17'd65621: data = 8'hef;
      17'd65622: data = 8'hed;
      17'd65623: data = 8'hed;
      17'd65624: data = 8'hf2;
      17'd65625: data = 8'hf5;
      17'd65626: data = 8'hfa;
      17'd65627: data = 8'hfa;
      17'd65628: data = 8'hf9;
      17'd65629: data = 8'hf6;
      17'd65630: data = 8'hfa;
      17'd65631: data = 8'hfe;
      17'd65632: data = 8'h01;
      17'd65633: data = 8'h04;
      17'd65634: data = 8'hfe;
      17'd65635: data = 8'hfa;
      17'd65636: data = 8'hf9;
      17'd65637: data = 8'hf9;
      17'd65638: data = 8'hfe;
      17'd65639: data = 8'h04;
      17'd65640: data = 8'h0a;
      17'd65641: data = 8'h06;
      17'd65642: data = 8'h06;
      17'd65643: data = 8'h05;
      17'd65644: data = 8'h02;
      17'd65645: data = 8'h05;
      17'd65646: data = 8'h0a;
      17'd65647: data = 8'h09;
      17'd65648: data = 8'h09;
      17'd65649: data = 8'h0a;
      17'd65650: data = 8'h05;
      17'd65651: data = 8'h05;
      17'd65652: data = 8'h09;
      17'd65653: data = 8'h0a;
      17'd65654: data = 8'h0c;
      17'd65655: data = 8'h0c;
      17'd65656: data = 8'h0c;
      17'd65657: data = 8'h0a;
      17'd65658: data = 8'h09;
      17'd65659: data = 8'h06;
      17'd65660: data = 8'h05;
      17'd65661: data = 8'h0c;
      17'd65662: data = 8'h0a;
      17'd65663: data = 8'h0a;
      17'd65664: data = 8'h0d;
      17'd65665: data = 8'h0c;
      17'd65666: data = 8'h0c;
      17'd65667: data = 8'h0a;
      17'd65668: data = 8'h09;
      17'd65669: data = 8'h04;
      17'd65670: data = 8'h02;
      17'd65671: data = 8'h09;
      17'd65672: data = 8'h0a;
      17'd65673: data = 8'h0a;
      17'd65674: data = 8'h0c;
      17'd65675: data = 8'h09;
      17'd65676: data = 8'h05;
      17'd65677: data = 8'h01;
      17'd65678: data = 8'hfe;
      17'd65679: data = 8'h00;
      17'd65680: data = 8'h00;
      17'd65681: data = 8'h01;
      17'd65682: data = 8'h02;
      17'd65683: data = 8'h00;
      17'd65684: data = 8'h00;
      17'd65685: data = 8'hfe;
      17'd65686: data = 8'hfd;
      17'd65687: data = 8'hfc;
      17'd65688: data = 8'hf9;
      17'd65689: data = 8'hf9;
      17'd65690: data = 8'hf6;
      17'd65691: data = 8'hf4;
      17'd65692: data = 8'hf6;
      17'd65693: data = 8'hfa;
      17'd65694: data = 8'hfc;
      17'd65695: data = 8'hf6;
      17'd65696: data = 8'hf4;
      17'd65697: data = 8'hf4;
      17'd65698: data = 8'hef;
      17'd65699: data = 8'hf1;
      17'd65700: data = 8'hf6;
      17'd65701: data = 8'hfa;
      17'd65702: data = 8'hfc;
      17'd65703: data = 8'hf9;
      17'd65704: data = 8'hf6;
      17'd65705: data = 8'hf2;
      17'd65706: data = 8'hed;
      17'd65707: data = 8'hef;
      17'd65708: data = 8'hf4;
      17'd65709: data = 8'hf4;
      17'd65710: data = 8'hf5;
      17'd65711: data = 8'hf4;
      17'd65712: data = 8'hf1;
      17'd65713: data = 8'hf4;
      17'd65714: data = 8'hf4;
      17'd65715: data = 8'hf4;
      17'd65716: data = 8'hf2;
      17'd65717: data = 8'hef;
      17'd65718: data = 8'hf6;
      17'd65719: data = 8'hf9;
      17'd65720: data = 8'hf9;
      17'd65721: data = 8'hfa;
      17'd65722: data = 8'hf9;
      17'd65723: data = 8'hf4;
      17'd65724: data = 8'hf2;
      17'd65725: data = 8'hf2;
      17'd65726: data = 8'hf2;
      17'd65727: data = 8'hf2;
      17'd65728: data = 8'hf1;
      17'd65729: data = 8'hfa;
      17'd65730: data = 8'h04;
      17'd65731: data = 8'h05;
      17'd65732: data = 8'h04;
      17'd65733: data = 8'h00;
      17'd65734: data = 8'hfe;
      17'd65735: data = 8'hfc;
      17'd65736: data = 8'hfc;
      17'd65737: data = 8'h02;
      17'd65738: data = 8'h05;
      17'd65739: data = 8'h02;
      17'd65740: data = 8'h04;
      17'd65741: data = 8'h0a;
      17'd65742: data = 8'h0c;
      17'd65743: data = 8'h04;
      17'd65744: data = 8'h01;
      17'd65745: data = 8'h05;
      17'd65746: data = 8'hfe;
      17'd65747: data = 8'h06;
      17'd65748: data = 8'h13;
      17'd65749: data = 8'h0e;
      17'd65750: data = 8'h0e;
      17'd65751: data = 8'h0e;
      17'd65752: data = 8'h0c;
      17'd65753: data = 8'h11;
      17'd65754: data = 8'h0c;
      17'd65755: data = 8'h0c;
      17'd65756: data = 8'h06;
      17'd65757: data = 8'h02;
      17'd65758: data = 8'h09;
      17'd65759: data = 8'h01;
      17'd65760: data = 8'h06;
      17'd65761: data = 8'h12;
      17'd65762: data = 8'h11;
      17'd65763: data = 8'h1b;
      17'd65764: data = 8'h19;
      17'd65765: data = 8'h0a;
      17'd65766: data = 8'h04;
      17'd65767: data = 8'h00;
      17'd65768: data = 8'h01;
      17'd65769: data = 8'h00;
      17'd65770: data = 8'h09;
      17'd65771: data = 8'h11;
      17'd65772: data = 8'h13;
      17'd65773: data = 8'h0d;
      17'd65774: data = 8'h01;
      17'd65775: data = 8'h01;
      17'd65776: data = 8'hfe;
      17'd65777: data = 8'hfa;
      17'd65778: data = 8'h00;
      17'd65779: data = 8'h04;
      17'd65780: data = 8'h02;
      17'd65781: data = 8'h01;
      17'd65782: data = 8'h05;
      17'd65783: data = 8'h01;
      17'd65784: data = 8'hfd;
      17'd65785: data = 8'h00;
      17'd65786: data = 8'hfd;
      17'd65787: data = 8'hf9;
      17'd65788: data = 8'hf2;
      17'd65789: data = 8'hfc;
      17'd65790: data = 8'hfc;
      17'd65791: data = 8'h00;
      17'd65792: data = 8'h06;
      17'd65793: data = 8'hfc;
      17'd65794: data = 8'h02;
      17'd65795: data = 8'h00;
      17'd65796: data = 8'hf2;
      17'd65797: data = 8'hfc;
      17'd65798: data = 8'hfd;
      17'd65799: data = 8'hfe;
      17'd65800: data = 8'h02;
      17'd65801: data = 8'h06;
      17'd65802: data = 8'hfd;
      17'd65803: data = 8'hf2;
      17'd65804: data = 8'hf4;
      17'd65805: data = 8'hf4;
      17'd65806: data = 8'h00;
      17'd65807: data = 8'h05;
      17'd65808: data = 8'h06;
      17'd65809: data = 8'h02;
      17'd65810: data = 8'h02;
      17'd65811: data = 8'h01;
      17'd65812: data = 8'hf4;
      17'd65813: data = 8'h00;
      17'd65814: data = 8'h04;
      17'd65815: data = 8'hfc;
      17'd65816: data = 8'hfa;
      17'd65817: data = 8'hf6;
      17'd65818: data = 8'hf1;
      17'd65819: data = 8'hf6;
      17'd65820: data = 8'h09;
      17'd65821: data = 8'h0a;
      17'd65822: data = 8'h0d;
      17'd65823: data = 8'h1a;
      17'd65824: data = 8'h05;
      17'd65825: data = 8'hf4;
      17'd65826: data = 8'hfc;
      17'd65827: data = 8'hfa;
      17'd65828: data = 8'hf9;
      17'd65829: data = 8'h0a;
      17'd65830: data = 8'h12;
      17'd65831: data = 8'h01;
      17'd65832: data = 8'hfd;
      17'd65833: data = 8'hfd;
      17'd65834: data = 8'hfd;
      17'd65835: data = 8'h06;
      17'd65836: data = 8'h16;
      17'd65837: data = 8'h15;
      17'd65838: data = 8'h05;
      17'd65839: data = 8'h01;
      17'd65840: data = 8'hf6;
      17'd65841: data = 8'hf5;
      17'd65842: data = 8'h04;
      17'd65843: data = 8'h11;
      17'd65844: data = 8'h13;
      17'd65845: data = 8'h12;
      17'd65846: data = 8'h04;
      17'd65847: data = 8'hf1;
      17'd65848: data = 8'hf4;
      17'd65849: data = 8'hfc;
      17'd65850: data = 8'h00;
      17'd65851: data = 8'h09;
      17'd65852: data = 8'h09;
      17'd65853: data = 8'hfd;
      17'd65854: data = 8'hf1;
      17'd65855: data = 8'hef;
      17'd65856: data = 8'hf4;
      17'd65857: data = 8'hfe;
      17'd65858: data = 8'h05;
      17'd65859: data = 8'h01;
      17'd65860: data = 8'hf4;
      17'd65861: data = 8'heb;
      17'd65862: data = 8'he3;
      17'd65863: data = 8'he2;
      17'd65864: data = 8'hec;
      17'd65865: data = 8'hf5;
      17'd65866: data = 8'hf6;
      17'd65867: data = 8'hf6;
      17'd65868: data = 8'hf1;
      17'd65869: data = 8'he7;
      17'd65870: data = 8'he7;
      17'd65871: data = 8'hf2;
      17'd65872: data = 8'hf2;
      17'd65873: data = 8'hf2;
      17'd65874: data = 8'hf2;
      17'd65875: data = 8'he5;
      17'd65876: data = 8'hde;
      17'd65877: data = 8'he2;
      17'd65878: data = 8'he9;
      17'd65879: data = 8'hf4;
      17'd65880: data = 8'hfc;
      17'd65881: data = 8'hfc;
      17'd65882: data = 8'hf6;
      17'd65883: data = 8'hf4;
      17'd65884: data = 8'hf4;
      17'd65885: data = 8'hf4;
      17'd65886: data = 8'hf5;
      17'd65887: data = 8'hfa;
      17'd65888: data = 8'hfa;
      17'd65889: data = 8'hf6;
      17'd65890: data = 8'hf6;
      17'd65891: data = 8'hf6;
      17'd65892: data = 8'hfc;
      17'd65893: data = 8'h04;
      17'd65894: data = 8'h06;
      17'd65895: data = 8'h05;
      17'd65896: data = 8'h04;
      17'd65897: data = 8'h02;
      17'd65898: data = 8'hfe;
      17'd65899: data = 8'h01;
      17'd65900: data = 8'h06;
      17'd65901: data = 8'h09;
      17'd65902: data = 8'h0d;
      17'd65903: data = 8'h0d;
      17'd65904: data = 8'h0c;
      17'd65905: data = 8'h0e;
      17'd65906: data = 8'h09;
      17'd65907: data = 8'h06;
      17'd65908: data = 8'h09;
      17'd65909: data = 8'h09;
      17'd65910: data = 8'h09;
      17'd65911: data = 8'h0a;
      17'd65912: data = 8'h0d;
      17'd65913: data = 8'h0e;
      17'd65914: data = 8'h0e;
      17'd65915: data = 8'h11;
      17'd65916: data = 8'h12;
      17'd65917: data = 8'h0a;
      17'd65918: data = 8'h0d;
      17'd65919: data = 8'h12;
      17'd65920: data = 8'h09;
      17'd65921: data = 8'h06;
      17'd65922: data = 8'h05;
      17'd65923: data = 8'h01;
      17'd65924: data = 8'h01;
      17'd65925: data = 8'h09;
      17'd65926: data = 8'h0a;
      17'd65927: data = 8'h0a;
      17'd65928: data = 8'h11;
      17'd65929: data = 8'h0d;
      17'd65930: data = 8'h04;
      17'd65931: data = 8'h04;
      17'd65932: data = 8'hfd;
      17'd65933: data = 8'hf9;
      17'd65934: data = 8'h01;
      17'd65935: data = 8'hfc;
      17'd65936: data = 8'hf6;
      17'd65937: data = 8'h02;
      17'd65938: data = 8'h00;
      17'd65939: data = 8'hfd;
      17'd65940: data = 8'hfd;
      17'd65941: data = 8'hfd;
      17'd65942: data = 8'hf6;
      17'd65943: data = 8'hf4;
      17'd65944: data = 8'hf2;
      17'd65945: data = 8'hef;
      17'd65946: data = 8'hf4;
      17'd65947: data = 8'hf6;
      17'd65948: data = 8'hf9;
      17'd65949: data = 8'hf5;
      17'd65950: data = 8'hf5;
      17'd65951: data = 8'hf1;
      17'd65952: data = 8'heb;
      17'd65953: data = 8'heb;
      17'd65954: data = 8'heb;
      17'd65955: data = 8'he7;
      17'd65956: data = 8'heb;
      17'd65957: data = 8'hed;
      17'd65958: data = 8'hed;
      17'd65959: data = 8'hf2;
      17'd65960: data = 8'hf5;
      17'd65961: data = 8'hed;
      17'd65962: data = 8'hef;
      17'd65963: data = 8'hf5;
      17'd65964: data = 8'hef;
      17'd65965: data = 8'hec;
      17'd65966: data = 8'heb;
      17'd65967: data = 8'he9;
      17'd65968: data = 8'hec;
      17'd65969: data = 8'hef;
      17'd65970: data = 8'hef;
      17'd65971: data = 8'hf4;
      17'd65972: data = 8'hf4;
      17'd65973: data = 8'hf2;
      17'd65974: data = 8'hf6;
      17'd65975: data = 8'hf2;
      17'd65976: data = 8'hf5;
      17'd65977: data = 8'hfa;
      17'd65978: data = 8'hf6;
      17'd65979: data = 8'hf4;
      17'd65980: data = 8'hf5;
      17'd65981: data = 8'hf9;
      17'd65982: data = 8'hfa;
      17'd65983: data = 8'hfc;
      17'd65984: data = 8'h00;
      17'd65985: data = 8'h00;
      17'd65986: data = 8'hfe;
      17'd65987: data = 8'h02;
      17'd65988: data = 8'h04;
      17'd65989: data = 8'h04;
      17'd65990: data = 8'h05;
      17'd65991: data = 8'h05;
      17'd65992: data = 8'h05;
      17'd65993: data = 8'h09;
      17'd65994: data = 8'h0e;
      17'd65995: data = 8'h0d;
      17'd65996: data = 8'h0c;
      17'd65997: data = 8'h0e;
      17'd65998: data = 8'h12;
      17'd65999: data = 8'h12;
      17'd66000: data = 8'h13;
      17'd66001: data = 8'h11;
      17'd66002: data = 8'h0c;
      17'd66003: data = 8'h0c;
      17'd66004: data = 8'h0e;
      17'd66005: data = 8'h12;
      17'd66006: data = 8'h16;
      17'd66007: data = 8'h1c;
      17'd66008: data = 8'h1b;
      17'd66009: data = 8'h13;
      17'd66010: data = 8'h13;
      17'd66011: data = 8'h13;
      17'd66012: data = 8'h11;
      17'd66013: data = 8'h11;
      17'd66014: data = 8'h11;
      17'd66015: data = 8'h0c;
      17'd66016: data = 8'h0c;
      17'd66017: data = 8'h13;
      17'd66018: data = 8'h0e;
      17'd66019: data = 8'h0e;
      17'd66020: data = 8'h15;
      17'd66021: data = 8'h15;
      17'd66022: data = 8'h12;
      17'd66023: data = 8'h13;
      17'd66024: data = 8'h0a;
      17'd66025: data = 8'h00;
      17'd66026: data = 8'h01;
      17'd66027: data = 8'hfa;
      17'd66028: data = 8'hfc;
      17'd66029: data = 8'h05;
      17'd66030: data = 8'h09;
      17'd66031: data = 8'h11;
      17'd66032: data = 8'h0e;
      17'd66033: data = 8'h09;
      17'd66034: data = 8'h02;
      17'd66035: data = 8'h05;
      17'd66036: data = 8'h00;
      17'd66037: data = 8'hf1;
      17'd66038: data = 8'hfd;
      17'd66039: data = 8'hfd;
      17'd66040: data = 8'hf2;
      17'd66041: data = 8'h00;
      17'd66042: data = 8'h0d;
      17'd66043: data = 8'h01;
      17'd66044: data = 8'h01;
      17'd66045: data = 8'h06;
      17'd66046: data = 8'hf4;
      17'd66047: data = 8'hf4;
      17'd66048: data = 8'hfa;
      17'd66049: data = 8'hf4;
      17'd66050: data = 8'hfd;
      17'd66051: data = 8'h0c;
      17'd66052: data = 8'h02;
      17'd66053: data = 8'h06;
      17'd66054: data = 8'h13;
      17'd66055: data = 8'h01;
      17'd66056: data = 8'h02;
      17'd66057: data = 8'h06;
      17'd66058: data = 8'hf5;
      17'd66059: data = 8'hfa;
      17'd66060: data = 8'hfe;
      17'd66061: data = 8'hfd;
      17'd66062: data = 8'hfa;
      17'd66063: data = 8'hfe;
      17'd66064: data = 8'h05;
      17'd66065: data = 8'h00;
      17'd66066: data = 8'h11;
      17'd66067: data = 8'h19;
      17'd66068: data = 8'h06;
      17'd66069: data = 8'h09;
      17'd66070: data = 8'h02;
      17'd66071: data = 8'hf2;
      17'd66072: data = 8'hf9;
      17'd66073: data = 8'h02;
      17'd66074: data = 8'hfe;
      17'd66075: data = 8'h0c;
      17'd66076: data = 8'h1a;
      17'd66077: data = 8'h0c;
      17'd66078: data = 8'h0c;
      17'd66079: data = 8'h0e;
      17'd66080: data = 8'h02;
      17'd66081: data = 8'h04;
      17'd66082: data = 8'h0d;
      17'd66083: data = 8'h02;
      17'd66084: data = 8'h05;
      17'd66085: data = 8'h0c;
      17'd66086: data = 8'h02;
      17'd66087: data = 8'h05;
      17'd66088: data = 8'h12;
      17'd66089: data = 8'h15;
      17'd66090: data = 8'h11;
      17'd66091: data = 8'h13;
      17'd66092: data = 8'h0a;
      17'd66093: data = 8'hfc;
      17'd66094: data = 8'hfe;
      17'd66095: data = 8'h01;
      17'd66096: data = 8'h02;
      17'd66097: data = 8'h0d;
      17'd66098: data = 8'h0e;
      17'd66099: data = 8'h04;
      17'd66100: data = 8'h02;
      17'd66101: data = 8'h04;
      17'd66102: data = 8'h01;
      17'd66103: data = 8'h01;
      17'd66104: data = 8'h02;
      17'd66105: data = 8'hfe;
      17'd66106: data = 8'hf9;
      17'd66107: data = 8'hf2;
      17'd66108: data = 8'heb;
      17'd66109: data = 8'heb;
      17'd66110: data = 8'hf2;
      17'd66111: data = 8'hf6;
      17'd66112: data = 8'hf9;
      17'd66113: data = 8'hf6;
      17'd66114: data = 8'hf2;
      17'd66115: data = 8'he9;
      17'd66116: data = 8'he5;
      17'd66117: data = 8'he5;
      17'd66118: data = 8'he3;
      17'd66119: data = 8'he5;
      17'd66120: data = 8'he4;
      17'd66121: data = 8'he0;
      17'd66122: data = 8'he2;
      17'd66123: data = 8'he4;
      17'd66124: data = 8'he3;
      17'd66125: data = 8'heb;
      17'd66126: data = 8'hf1;
      17'd66127: data = 8'hec;
      17'd66128: data = 8'he9;
      17'd66129: data = 8'he2;
      17'd66130: data = 8'hdb;
      17'd66131: data = 8'hdb;
      17'd66132: data = 8'he3;
      17'd66133: data = 8'hec;
      17'd66134: data = 8'hf2;
      17'd66135: data = 8'hf9;
      17'd66136: data = 8'hfa;
      17'd66137: data = 8'hf6;
      17'd66138: data = 8'hf9;
      17'd66139: data = 8'hf6;
      17'd66140: data = 8'hf6;
      17'd66141: data = 8'hf6;
      17'd66142: data = 8'hfa;
      17'd66143: data = 8'hf9;
      17'd66144: data = 8'hfa;
      17'd66145: data = 8'h01;
      17'd66146: data = 8'h05;
      17'd66147: data = 8'h0a;
      17'd66148: data = 8'h0e;
      17'd66149: data = 8'h0e;
      17'd66150: data = 8'h0e;
      17'd66151: data = 8'h11;
      17'd66152: data = 8'h0c;
      17'd66153: data = 8'h0c;
      17'd66154: data = 8'h0e;
      17'd66155: data = 8'h11;
      17'd66156: data = 8'h11;
      17'd66157: data = 8'h15;
      17'd66158: data = 8'h1a;
      17'd66159: data = 8'h19;
      17'd66160: data = 8'h1a;
      17'd66161: data = 8'h1b;
      17'd66162: data = 8'h1a;
      17'd66163: data = 8'h1a;
      17'd66164: data = 8'h15;
      17'd66165: data = 8'h13;
      17'd66166: data = 8'h0e;
      17'd66167: data = 8'h0c;
      17'd66168: data = 8'h0e;
      17'd66169: data = 8'h0e;
      17'd66170: data = 8'h19;
      17'd66171: data = 8'h1a;
      17'd66172: data = 8'h13;
      17'd66173: data = 8'h11;
      17'd66174: data = 8'h0d;
      17'd66175: data = 8'h01;
      17'd66176: data = 8'h00;
      17'd66177: data = 8'h06;
      17'd66178: data = 8'h02;
      17'd66179: data = 8'h02;
      17'd66180: data = 8'h09;
      17'd66181: data = 8'hfe;
      17'd66182: data = 8'hf2;
      17'd66183: data = 8'hfc;
      17'd66184: data = 8'hfc;
      17'd66185: data = 8'hfa;
      17'd66186: data = 8'h02;
      17'd66187: data = 8'h00;
      17'd66188: data = 8'hfa;
      17'd66189: data = 8'hf5;
      17'd66190: data = 8'heb;
      17'd66191: data = 8'he5;
      17'd66192: data = 8'heb;
      17'd66193: data = 8'hec;
      17'd66194: data = 8'he7;
      17'd66195: data = 8'heb;
      17'd66196: data = 8'he9;
      17'd66197: data = 8'he4;
      17'd66198: data = 8'hec;
      17'd66199: data = 8'hec;
      17'd66200: data = 8'hec;
      17'd66201: data = 8'hec;
      17'd66202: data = 8'he4;
      17'd66203: data = 8'he0;
      17'd66204: data = 8'hd3;
      17'd66205: data = 8'hd5;
      17'd66206: data = 8'he0;
      17'd66207: data = 8'he2;
      17'd66208: data = 8'heb;
      17'd66209: data = 8'hed;
      17'd66210: data = 8'he7;
      17'd66211: data = 8'he0;
      17'd66212: data = 8'he0;
      17'd66213: data = 8'hde;
      17'd66214: data = 8'he0;
      17'd66215: data = 8'he5;
      17'd66216: data = 8'he2;
      17'd66217: data = 8'he4;
      17'd66218: data = 8'he9;
      17'd66219: data = 8'he7;
      17'd66220: data = 8'hed;
      17'd66221: data = 8'hf2;
      17'd66222: data = 8'hf1;
      17'd66223: data = 8'hf4;
      17'd66224: data = 8'hf2;
      17'd66225: data = 8'heb;
      17'd66226: data = 8'he7;
      17'd66227: data = 8'hef;
      17'd66228: data = 8'hf4;
      17'd66229: data = 8'hfc;
      17'd66230: data = 8'h01;
      17'd66231: data = 8'h00;
      17'd66232: data = 8'h02;
      17'd66233: data = 8'hfe;
      17'd66234: data = 8'hfd;
      17'd66235: data = 8'h01;
      17'd66236: data = 8'h05;
      17'd66237: data = 8'h05;
      17'd66238: data = 8'h09;
      17'd66239: data = 8'h0a;
      17'd66240: data = 8'h0a;
      17'd66241: data = 8'h0a;
      17'd66242: data = 8'h0c;
      17'd66243: data = 8'h11;
      17'd66244: data = 8'h12;
      17'd66245: data = 8'h13;
      17'd66246: data = 8'h15;
      17'd66247: data = 8'h12;
      17'd66248: data = 8'h15;
      17'd66249: data = 8'h15;
      17'd66250: data = 8'h16;
      17'd66251: data = 8'h1a;
      17'd66252: data = 8'h15;
      17'd66253: data = 8'h15;
      17'd66254: data = 8'h12;
      17'd66255: data = 8'h0e;
      17'd66256: data = 8'h13;
      17'd66257: data = 8'h1b;
      17'd66258: data = 8'h1b;
      17'd66259: data = 8'h1e;
      17'd66260: data = 8'h1a;
      17'd66261: data = 8'h15;
      17'd66262: data = 8'h11;
      17'd66263: data = 8'h11;
      17'd66264: data = 8'h0d;
      17'd66265: data = 8'h09;
      17'd66266: data = 8'h0e;
      17'd66267: data = 8'h0c;
      17'd66268: data = 8'h11;
      17'd66269: data = 8'h19;
      17'd66270: data = 8'h11;
      17'd66271: data = 8'h0e;
      17'd66272: data = 8'h11;
      17'd66273: data = 8'h06;
      17'd66274: data = 8'h02;
      17'd66275: data = 8'h02;
      17'd66276: data = 8'h00;
      17'd66277: data = 8'h02;
      17'd66278: data = 8'h06;
      17'd66279: data = 8'h06;
      17'd66280: data = 8'h0a;
      17'd66281: data = 8'h0c;
      17'd66282: data = 8'h05;
      17'd66283: data = 8'hfe;
      17'd66284: data = 8'hfd;
      17'd66285: data = 8'hf9;
      17'd66286: data = 8'hfc;
      17'd66287: data = 8'h00;
      17'd66288: data = 8'h04;
      17'd66289: data = 8'h01;
      17'd66290: data = 8'hfc;
      17'd66291: data = 8'h05;
      17'd66292: data = 8'hf9;
      17'd66293: data = 8'hf6;
      17'd66294: data = 8'h01;
      17'd66295: data = 8'h04;
      17'd66296: data = 8'h00;
      17'd66297: data = 8'hfc;
      17'd66298: data = 8'h0c;
      17'd66299: data = 8'h00;
      17'd66300: data = 8'h05;
      17'd66301: data = 8'h09;
      17'd66302: data = 8'hfe;
      17'd66303: data = 8'h05;
      17'd66304: data = 8'hfa;
      17'd66305: data = 8'hf5;
      17'd66306: data = 8'h05;
      17'd66307: data = 8'h06;
      17'd66308: data = 8'h01;
      17'd66309: data = 8'h0a;
      17'd66310: data = 8'h0a;
      17'd66311: data = 8'hfd;
      17'd66312: data = 8'hf5;
      17'd66313: data = 8'hfa;
      17'd66314: data = 8'h01;
      17'd66315: data = 8'h05;
      17'd66316: data = 8'h1b;
      17'd66317: data = 8'h15;
      17'd66318: data = 8'h0d;
      17'd66319: data = 8'h0c;
      17'd66320: data = 8'hf9;
      17'd66321: data = 8'hfd;
      17'd66322: data = 8'hf9;
      17'd66323: data = 8'hfc;
      17'd66324: data = 8'h0e;
      17'd66325: data = 8'h12;
      17'd66326: data = 8'h11;
      17'd66327: data = 8'h12;
      17'd66328: data = 8'h0e;
      17'd66329: data = 8'h12;
      17'd66330: data = 8'h13;
      17'd66331: data = 8'h0c;
      17'd66332: data = 8'h06;
      17'd66333: data = 8'h00;
      17'd66334: data = 8'hf5;
      17'd66335: data = 8'hfa;
      17'd66336: data = 8'h09;
      17'd66337: data = 8'h15;
      17'd66338: data = 8'h1c;
      17'd66339: data = 8'h1f;
      17'd66340: data = 8'h12;
      17'd66341: data = 8'h04;
      17'd66342: data = 8'hfe;
      17'd66343: data = 8'hf5;
      17'd66344: data = 8'hfd;
      17'd66345: data = 8'h00;
      17'd66346: data = 8'h01;
      17'd66347: data = 8'h05;
      17'd66348: data = 8'hfa;
      17'd66349: data = 8'hf9;
      17'd66350: data = 8'h04;
      17'd66351: data = 8'h01;
      17'd66352: data = 8'hfd;
      17'd66353: data = 8'h00;
      17'd66354: data = 8'hf4;
      17'd66355: data = 8'he9;
      17'd66356: data = 8'he3;
      17'd66357: data = 8'hdb;
      17'd66358: data = 8'he4;
      17'd66359: data = 8'hec;
      17'd66360: data = 8'hef;
      17'd66361: data = 8'hec;
      17'd66362: data = 8'he4;
      17'd66363: data = 8'hda;
      17'd66364: data = 8'hd5;
      17'd66365: data = 8'hda;
      17'd66366: data = 8'hda;
      17'd66367: data = 8'he0;
      17'd66368: data = 8'he2;
      17'd66369: data = 8'hdb;
      17'd66370: data = 8'hd5;
      17'd66371: data = 8'hd3;
      17'd66372: data = 8'hd3;
      17'd66373: data = 8'hd8;
      17'd66374: data = 8'hde;
      17'd66375: data = 8'hde;
      17'd66376: data = 8'he4;
      17'd66377: data = 8'he0;
      17'd66378: data = 8'hda;
      17'd66379: data = 8'he4;
      17'd66380: data = 8'he7;
      17'd66381: data = 8'hec;
      17'd66382: data = 8'hf1;
      17'd66383: data = 8'hed;
      17'd66384: data = 8'hec;
      17'd66385: data = 8'hef;
      17'd66386: data = 8'hf2;
      17'd66387: data = 8'hf9;
      17'd66388: data = 8'h02;
      17'd66389: data = 8'h09;
      17'd66390: data = 8'h0e;
      17'd66391: data = 8'h0a;
      17'd66392: data = 8'h04;
      17'd66393: data = 8'h06;
      17'd66394: data = 8'h06;
      17'd66395: data = 8'h09;
      17'd66396: data = 8'h11;
      17'd66397: data = 8'h19;
      17'd66398: data = 8'h1c;
      17'd66399: data = 8'h1f;
      17'd66400: data = 8'h22;
      17'd66401: data = 8'h1e;
      17'd66402: data = 8'h1e;
      17'd66403: data = 8'h1e;
      17'd66404: data = 8'h1a;
      17'd66405: data = 8'h1b;
      17'd66406: data = 8'h1a;
      17'd66407: data = 8'h16;
      17'd66408: data = 8'h1a;
      17'd66409: data = 8'h1c;
      17'd66410: data = 8'h22;
      17'd66411: data = 8'h29;
      17'd66412: data = 8'h22;
      17'd66413: data = 8'h19;
      17'd66414: data = 8'h1a;
      17'd66415: data = 8'h0e;
      17'd66416: data = 8'h0a;
      17'd66417: data = 8'h0d;
      17'd66418: data = 8'h0e;
      17'd66419: data = 8'h11;
      17'd66420: data = 8'h0d;
      17'd66421: data = 8'h0e;
      17'd66422: data = 8'h0a;
      17'd66423: data = 8'h05;
      17'd66424: data = 8'h04;
      17'd66425: data = 8'h01;
      17'd66426: data = 8'h01;
      17'd66427: data = 8'hf4;
      17'd66428: data = 8'hef;
      17'd66429: data = 8'hf2;
      17'd66430: data = 8'hed;
      17'd66431: data = 8'hf5;
      17'd66432: data = 8'hf6;
      17'd66433: data = 8'hf1;
      17'd66434: data = 8'hed;
      17'd66435: data = 8'he7;
      17'd66436: data = 8'he3;
      17'd66437: data = 8'he2;
      17'd66438: data = 8'he0;
      17'd66439: data = 8'he0;
      17'd66440: data = 8'he3;
      17'd66441: data = 8'he0;
      17'd66442: data = 8'hdb;
      17'd66443: data = 8'he0;
      17'd66444: data = 8'hdc;
      17'd66445: data = 8'hdc;
      17'd66446: data = 8'hdc;
      17'd66447: data = 8'hda;
      17'd66448: data = 8'hda;
      17'd66449: data = 8'hda;
      17'd66450: data = 8'hda;
      17'd66451: data = 8'hdb;
      17'd66452: data = 8'hde;
      17'd66453: data = 8'hdc;
      17'd66454: data = 8'hdb;
      17'd66455: data = 8'hdc;
      17'd66456: data = 8'hd8;
      17'd66457: data = 8'he0;
      17'd66458: data = 8'he4;
      17'd66459: data = 8'he2;
      17'd66460: data = 8'he9;
      17'd66461: data = 8'hed;
      17'd66462: data = 8'hec;
      17'd66463: data = 8'hec;
      17'd66464: data = 8'hec;
      17'd66465: data = 8'hed;
      17'd66466: data = 8'hed;
      17'd66467: data = 8'hef;
      17'd66468: data = 8'hf2;
      17'd66469: data = 8'hf9;
      17'd66470: data = 8'hfe;
      17'd66471: data = 8'h01;
      17'd66472: data = 8'h02;
      17'd66473: data = 8'h00;
      17'd66474: data = 8'h04;
      17'd66475: data = 8'h01;
      17'd66476: data = 8'h02;
      17'd66477: data = 8'h01;
      17'd66478: data = 8'h01;
      17'd66479: data = 8'h0a;
      17'd66480: data = 8'h0d;
      17'd66481: data = 8'h12;
      17'd66482: data = 8'h15;
      17'd66483: data = 8'h15;
      17'd66484: data = 8'h16;
      17'd66485: data = 8'h13;
      17'd66486: data = 8'h13;
      17'd66487: data = 8'h15;
      17'd66488: data = 8'h16;
      17'd66489: data = 8'h15;
      17'd66490: data = 8'h13;
      17'd66491: data = 8'h16;
      17'd66492: data = 8'h16;
      17'd66493: data = 8'h1a;
      17'd66494: data = 8'h1b;
      17'd66495: data = 8'h1c;
      17'd66496: data = 8'h1c;
      17'd66497: data = 8'h15;
      17'd66498: data = 8'h15;
      17'd66499: data = 8'h15;
      17'd66500: data = 8'h12;
      17'd66501: data = 8'h12;
      17'd66502: data = 8'h15;
      17'd66503: data = 8'h12;
      17'd66504: data = 8'h0e;
      17'd66505: data = 8'h12;
      17'd66506: data = 8'h06;
      17'd66507: data = 8'h09;
      17'd66508: data = 8'h13;
      17'd66509: data = 8'h09;
      17'd66510: data = 8'h0c;
      17'd66511: data = 8'h0d;
      17'd66512: data = 8'h04;
      17'd66513: data = 8'h0c;
      17'd66514: data = 8'h04;
      17'd66515: data = 8'h00;
      17'd66516: data = 8'h01;
      17'd66517: data = 8'h06;
      17'd66518: data = 8'hfe;
      17'd66519: data = 8'hfd;
      17'd66520: data = 8'h06;
      17'd66521: data = 8'hf9;
      17'd66522: data = 8'h04;
      17'd66523: data = 8'h02;
      17'd66524: data = 8'hfd;
      17'd66525: data = 8'h0a;
      17'd66526: data = 8'hfe;
      17'd66527: data = 8'hfd;
      17'd66528: data = 8'h04;
      17'd66529: data = 8'h04;
      17'd66530: data = 8'hfc;
      17'd66531: data = 8'h11;
      17'd66532: data = 8'h09;
      17'd66533: data = 8'hf9;
      17'd66534: data = 8'h12;
      17'd66535: data = 8'hfe;
      17'd66536: data = 8'hfd;
      17'd66537: data = 8'h11;
      17'd66538: data = 8'h05;
      17'd66539: data = 8'h0c;
      17'd66540: data = 8'h0a;
      17'd66541: data = 8'h06;
      17'd66542: data = 8'h0d;
      17'd66543: data = 8'h11;
      17'd66544: data = 8'h09;
      17'd66545: data = 8'h09;
      17'd66546: data = 8'h0e;
      17'd66547: data = 8'h02;
      17'd66548: data = 8'h00;
      17'd66549: data = 8'h11;
      17'd66550: data = 8'h0d;
      17'd66551: data = 8'h16;
      17'd66552: data = 8'h19;
      17'd66553: data = 8'h02;
      17'd66554: data = 8'h0a;
      17'd66555: data = 8'hf5;
      17'd66556: data = 8'he5;
      17'd66557: data = 8'h06;
      17'd66558: data = 8'h05;
      17'd66559: data = 8'h12;
      17'd66560: data = 8'h26;
      17'd66561: data = 8'h1b;
      17'd66562: data = 8'h15;
      17'd66563: data = 8'h12;
      17'd66564: data = 8'h05;
      17'd66565: data = 8'h00;
      17'd66566: data = 8'h0c;
      17'd66567: data = 8'h0a;
      17'd66568: data = 8'h05;
      17'd66569: data = 8'h11;
      17'd66570: data = 8'h05;
      17'd66571: data = 8'h09;
      17'd66572: data = 8'h24;
      17'd66573: data = 8'h1f;
      17'd66574: data = 8'h22;
      17'd66575: data = 8'h26;
      17'd66576: data = 8'h0d;
      17'd66577: data = 8'h01;
      17'd66578: data = 8'hfe;
      17'd66579: data = 8'hfd;
      17'd66580: data = 8'h13;
      17'd66581: data = 8'h1b;
      17'd66582: data = 8'h19;
      17'd66583: data = 8'h1a;
      17'd66584: data = 8'h0d;
      17'd66585: data = 8'h00;
      17'd66586: data = 8'h02;
      17'd66587: data = 8'h0a;
      17'd66588: data = 8'h0a;
      17'd66589: data = 8'h0e;
      17'd66590: data = 8'h0d;
      17'd66591: data = 8'hfc;
      17'd66592: data = 8'hf5;
      17'd66593: data = 8'hf5;
      17'd66594: data = 8'hf6;
      17'd66595: data = 8'hfd;
      17'd66596: data = 8'hf4;
      17'd66597: data = 8'hec;
      17'd66598: data = 8'heb;
      17'd66599: data = 8'hdb;
      17'd66600: data = 8'hdc;
      17'd66601: data = 8'he9;
      17'd66602: data = 8'he9;
      17'd66603: data = 8'hef;
      17'd66604: data = 8'he9;
      17'd66605: data = 8'hdb;
      17'd66606: data = 8'hd2;
      17'd66607: data = 8'hc9;
      17'd66608: data = 8'hc6;
      17'd66609: data = 8'hce;
      17'd66610: data = 8'hd8;
      17'd66611: data = 8'hd8;
      17'd66612: data = 8'he0;
      17'd66613: data = 8'hde;
      17'd66614: data = 8'hd3;
      17'd66615: data = 8'hda;
      17'd66616: data = 8'hdb;
      17'd66617: data = 8'hda;
      17'd66618: data = 8'hdc;
      17'd66619: data = 8'hdc;
      17'd66620: data = 8'hdb;
      17'd66621: data = 8'hdc;
      17'd66622: data = 8'he3;
      17'd66623: data = 8'he9;
      17'd66624: data = 8'hfc;
      17'd66625: data = 8'hfe;
      17'd66626: data = 8'hfc;
      17'd66627: data = 8'hfc;
      17'd66628: data = 8'hfa;
      17'd66629: data = 8'hfc;
      17'd66630: data = 8'hfe;
      17'd66631: data = 8'h05;
      17'd66632: data = 8'h09;
      17'd66633: data = 8'h12;
      17'd66634: data = 8'h12;
      17'd66635: data = 8'h12;
      17'd66636: data = 8'h19;
      17'd66637: data = 8'h16;
      17'd66638: data = 8'h1a;
      17'd66639: data = 8'h1c;
      17'd66640: data = 8'h1a;
      17'd66641: data = 8'h1f;
      17'd66642: data = 8'h23;
      17'd66643: data = 8'h22;
      17'd66644: data = 8'h26;
      17'd66645: data = 8'h26;
      17'd66646: data = 8'h26;
      17'd66647: data = 8'h24;
      17'd66648: data = 8'h1e;
      17'd66649: data = 8'h1c;
      17'd66650: data = 8'h1b;
      17'd66651: data = 8'h1a;
      17'd66652: data = 8'h1a;
      17'd66653: data = 8'h1e;
      17'd66654: data = 8'h1f;
      17'd66655: data = 8'h1a;
      17'd66656: data = 8'h19;
      17'd66657: data = 8'h13;
      17'd66658: data = 8'h05;
      17'd66659: data = 8'h06;
      17'd66660: data = 8'h05;
      17'd66661: data = 8'hfd;
      17'd66662: data = 8'h02;
      17'd66663: data = 8'h01;
      17'd66664: data = 8'hfd;
      17'd66665: data = 8'hfd;
      17'd66666: data = 8'hf6;
      17'd66667: data = 8'hf5;
      17'd66668: data = 8'hf4;
      17'd66669: data = 8'hed;
      17'd66670: data = 8'he4;
      17'd66671: data = 8'he5;
      17'd66672: data = 8'hde;
      17'd66673: data = 8'hd5;
      17'd66674: data = 8'hde;
      17'd66675: data = 8'hdc;
      17'd66676: data = 8'hda;
      17'd66677: data = 8'hde;
      17'd66678: data = 8'hdc;
      17'd66679: data = 8'hd6;
      17'd66680: data = 8'hd8;
      17'd66681: data = 8'hda;
      17'd66682: data = 8'hd6;
      17'd66683: data = 8'hda;
      17'd66684: data = 8'hd6;
      17'd66685: data = 8'hd3;
      17'd66686: data = 8'hd3;
      17'd66687: data = 8'hce;
      17'd66688: data = 8'hd2;
      17'd66689: data = 8'hd6;
      17'd66690: data = 8'hda;
      17'd66691: data = 8'hdc;
      17'd66692: data = 8'he0;
      17'd66693: data = 8'he3;
      17'd66694: data = 8'he3;
      17'd66695: data = 8'he9;
      17'd66696: data = 8'he9;
      17'd66697: data = 8'heb;
      17'd66698: data = 8'hec;
      17'd66699: data = 8'he9;
      17'd66700: data = 8'hec;
      17'd66701: data = 8'hec;
      17'd66702: data = 8'hef;
      17'd66703: data = 8'hf5;
      17'd66704: data = 8'hf6;
      17'd66705: data = 8'hfe;
      17'd66706: data = 8'h02;
      17'd66707: data = 8'h04;
      17'd66708: data = 8'h04;
      17'd66709: data = 8'h0a;
      17'd66710: data = 8'h0a;
      17'd66711: data = 8'h09;
      17'd66712: data = 8'h0c;
      17'd66713: data = 8'h0a;
      17'd66714: data = 8'h0a;
      17'd66715: data = 8'h0e;
      17'd66716: data = 8'h0c;
      17'd66717: data = 8'h0d;
      17'd66718: data = 8'h0e;
      17'd66719: data = 8'h0e;
      17'd66720: data = 8'h13;
      17'd66721: data = 8'h16;
      17'd66722: data = 8'h16;
      17'd66723: data = 8'h19;
      17'd66724: data = 8'h1b;
      17'd66725: data = 8'h16;
      17'd66726: data = 8'h13;
      17'd66727: data = 8'h12;
      17'd66728: data = 8'h0a;
      17'd66729: data = 8'h0c;
      17'd66730: data = 8'h0e;
      17'd66731: data = 8'h0c;
      17'd66732: data = 8'h0e;
      17'd66733: data = 8'h12;
      17'd66734: data = 8'h0d;
      17'd66735: data = 8'h0a;
      17'd66736: data = 8'h0e;
      17'd66737: data = 8'h0d;
      17'd66738: data = 8'h0a;
      17'd66739: data = 8'h0c;
      17'd66740: data = 8'h06;
      17'd66741: data = 8'h02;
      17'd66742: data = 8'h01;
      17'd66743: data = 8'hfe;
      17'd66744: data = 8'hfe;
      17'd66745: data = 8'h00;
      17'd66746: data = 8'h01;
      17'd66747: data = 8'hfa;
      17'd66748: data = 8'h02;
      17'd66749: data = 8'h00;
      17'd66750: data = 8'hfe;
      17'd66751: data = 8'h09;
      17'd66752: data = 8'h01;
      17'd66753: data = 8'h02;
      17'd66754: data = 8'hfe;
      17'd66755: data = 8'hfe;
      17'd66756: data = 8'hf6;
      17'd66757: data = 8'hf9;
      17'd66758: data = 8'h01;
      17'd66759: data = 8'hf6;
      17'd66760: data = 8'h02;
      17'd66761: data = 8'h06;
      17'd66762: data = 8'h00;
      17'd66763: data = 8'h0c;
      17'd66764: data = 8'h09;
      17'd66765: data = 8'h09;
      17'd66766: data = 8'h0d;
      17'd66767: data = 8'h0d;
      17'd66768: data = 8'h09;
      17'd66769: data = 8'h0a;
      17'd66770: data = 8'h05;
      17'd66771: data = 8'h02;
      17'd66772: data = 8'h05;
      17'd66773: data = 8'h06;
      17'd66774: data = 8'h06;
      17'd66775: data = 8'h0d;
      17'd66776: data = 8'h1a;
      17'd66777: data = 8'h0c;
      17'd66778: data = 8'h15;
      17'd66779: data = 8'h1c;
      17'd66780: data = 8'h13;
      17'd66781: data = 8'h13;
      17'd66782: data = 8'h0d;
      17'd66783: data = 8'h11;
      17'd66784: data = 8'h09;
      17'd66785: data = 8'h09;
      17'd66786: data = 8'h0e;
      17'd66787: data = 8'h11;
      17'd66788: data = 8'h15;
      17'd66789: data = 8'h1b;
      17'd66790: data = 8'h1e;
      17'd66791: data = 8'h15;
      17'd66792: data = 8'h0a;
      17'd66793: data = 8'h00;
      17'd66794: data = 8'h01;
      17'd66795: data = 8'h00;
      17'd66796: data = 8'h00;
      17'd66797: data = 8'h12;
      17'd66798: data = 8'h16;
      17'd66799: data = 8'h16;
      17'd66800: data = 8'h11;
      17'd66801: data = 8'h0c;
      17'd66802: data = 8'h00;
      17'd66803: data = 8'hfd;
      17'd66804: data = 8'h02;
      17'd66805: data = 8'h04;
      17'd66806: data = 8'h0d;
      17'd66807: data = 8'h06;
      17'd66808: data = 8'h0c;
      17'd66809: data = 8'h0c;
      17'd66810: data = 8'h05;
      17'd66811: data = 8'h0c;
      17'd66812: data = 8'h0d;
      17'd66813: data = 8'h09;
      17'd66814: data = 8'h02;
      17'd66815: data = 8'h01;
      17'd66816: data = 8'h02;
      17'd66817: data = 8'h06;
      17'd66818: data = 8'h11;
      17'd66819: data = 8'h1e;
      17'd66820: data = 8'h24;
      17'd66821: data = 8'h15;
      17'd66822: data = 8'h04;
      17'd66823: data = 8'hfc;
      17'd66824: data = 8'hf5;
      17'd66825: data = 8'hf6;
      17'd66826: data = 8'h04;
      17'd66827: data = 8'h0c;
      17'd66828: data = 8'h12;
      17'd66829: data = 8'h15;
      17'd66830: data = 8'h09;
      17'd66831: data = 8'h09;
      17'd66832: data = 8'h09;
      17'd66833: data = 8'h05;
      17'd66834: data = 8'h06;
      17'd66835: data = 8'hfd;
      17'd66836: data = 8'hf2;
      17'd66837: data = 8'hf2;
      17'd66838: data = 8'hf2;
      17'd66839: data = 8'hf1;
      17'd66840: data = 8'hf6;
      17'd66841: data = 8'hfd;
      17'd66842: data = 8'hfc;
      17'd66843: data = 8'hf2;
      17'd66844: data = 8'he9;
      17'd66845: data = 8'he3;
      17'd66846: data = 8'he5;
      17'd66847: data = 8'he5;
      17'd66848: data = 8'he4;
      17'd66849: data = 8'hef;
      17'd66850: data = 8'hec;
      17'd66851: data = 8'he7;
      17'd66852: data = 8'he4;
      17'd66853: data = 8'hdc;
      17'd66854: data = 8'hda;
      17'd66855: data = 8'hda;
      17'd66856: data = 8'hdc;
      17'd66857: data = 8'hde;
      17'd66858: data = 8'he0;
      17'd66859: data = 8'he3;
      17'd66860: data = 8'heb;
      17'd66861: data = 8'hec;
      17'd66862: data = 8'hed;
      17'd66863: data = 8'hf1;
      17'd66864: data = 8'hf1;
      17'd66865: data = 8'hec;
      17'd66866: data = 8'he3;
      17'd66867: data = 8'he7;
      17'd66868: data = 8'he9;
      17'd66869: data = 8'hef;
      17'd66870: data = 8'hf5;
      17'd66871: data = 8'hfd;
      17'd66872: data = 8'h04;
      17'd66873: data = 8'h04;
      17'd66874: data = 8'h05;
      17'd66875: data = 8'h06;
      17'd66876: data = 8'h06;
      17'd66877: data = 8'h0a;
      17'd66878: data = 8'h0a;
      17'd66879: data = 8'h0a;
      17'd66880: data = 8'h0d;
      17'd66881: data = 8'h13;
      17'd66882: data = 8'h15;
      17'd66883: data = 8'h15;
      17'd66884: data = 8'h12;
      17'd66885: data = 8'h13;
      17'd66886: data = 8'h16;
      17'd66887: data = 8'h13;
      17'd66888: data = 8'h12;
      17'd66889: data = 8'h12;
      17'd66890: data = 8'h19;
      17'd66891: data = 8'h19;
      17'd66892: data = 8'h16;
      17'd66893: data = 8'h16;
      17'd66894: data = 8'h19;
      17'd66895: data = 8'h16;
      17'd66896: data = 8'h0e;
      17'd66897: data = 8'h09;
      17'd66898: data = 8'h01;
      17'd66899: data = 8'hfd;
      17'd66900: data = 8'hfc;
      17'd66901: data = 8'hfe;
      17'd66902: data = 8'h00;
      17'd66903: data = 8'h00;
      17'd66904: data = 8'h04;
      17'd66905: data = 8'hfe;
      17'd66906: data = 8'hfa;
      17'd66907: data = 8'hfa;
      17'd66908: data = 8'hf9;
      17'd66909: data = 8'hed;
      17'd66910: data = 8'he4;
      17'd66911: data = 8'he2;
      17'd66912: data = 8'he3;
      17'd66913: data = 8'he0;
      17'd66914: data = 8'he0;
      17'd66915: data = 8'he7;
      17'd66916: data = 8'he5;
      17'd66917: data = 8'he2;
      17'd66918: data = 8'hde;
      17'd66919: data = 8'hda;
      17'd66920: data = 8'hda;
      17'd66921: data = 8'hda;
      17'd66922: data = 8'hde;
      17'd66923: data = 8'he3;
      17'd66924: data = 8'he4;
      17'd66925: data = 8'he0;
      17'd66926: data = 8'hdb;
      17'd66927: data = 8'hdb;
      17'd66928: data = 8'hd6;
      17'd66929: data = 8'hda;
      17'd66930: data = 8'he0;
      17'd66931: data = 8'he0;
      17'd66932: data = 8'he5;
      17'd66933: data = 8'hec;
      17'd66934: data = 8'hed;
      17'd66935: data = 8'hf1;
      17'd66936: data = 8'hf6;
      17'd66937: data = 8'hf5;
      17'd66938: data = 8'hf2;
      17'd66939: data = 8'hed;
      17'd66940: data = 8'he7;
      17'd66941: data = 8'he9;
      17'd66942: data = 8'hed;
      17'd66943: data = 8'hf5;
      17'd66944: data = 8'hfd;
      17'd66945: data = 8'h00;
      17'd66946: data = 8'h02;
      17'd66947: data = 8'h00;
      17'd66948: data = 8'hfe;
      17'd66949: data = 8'h00;
      17'd66950: data = 8'h00;
      17'd66951: data = 8'h04;
      17'd66952: data = 8'h09;
      17'd66953: data = 8'h0e;
      17'd66954: data = 8'h0d;
      17'd66955: data = 8'h09;
      17'd66956: data = 8'h05;
      17'd66957: data = 8'h04;
      17'd66958: data = 8'h09;
      17'd66959: data = 8'h06;
      17'd66960: data = 8'h05;
      17'd66961: data = 8'h09;
      17'd66962: data = 8'h06;
      17'd66963: data = 8'h0a;
      17'd66964: data = 8'h11;
      17'd66965: data = 8'h12;
      17'd66966: data = 8'h11;
      17'd66967: data = 8'h0e;
      17'd66968: data = 8'h0a;
      17'd66969: data = 8'h05;
      17'd66970: data = 8'h00;
      17'd66971: data = 8'hfe;
      17'd66972: data = 8'h02;
      17'd66973: data = 8'h02;
      17'd66974: data = 8'h06;
      17'd66975: data = 8'h05;
      17'd66976: data = 8'h02;
      17'd66977: data = 8'h01;
      17'd66978: data = 8'h04;
      17'd66979: data = 8'h01;
      17'd66980: data = 8'h01;
      17'd66981: data = 8'h05;
      17'd66982: data = 8'h01;
      17'd66983: data = 8'h01;
      17'd66984: data = 8'h02;
      17'd66985: data = 8'h01;
      17'd66986: data = 8'h00;
      17'd66987: data = 8'h00;
      17'd66988: data = 8'hfc;
      17'd66989: data = 8'h00;
      17'd66990: data = 8'hfd;
      17'd66991: data = 8'hf9;
      17'd66992: data = 8'h02;
      17'd66993: data = 8'h00;
      17'd66994: data = 8'h05;
      17'd66995: data = 8'h0d;
      17'd66996: data = 8'h0a;
      17'd66997: data = 8'h09;
      17'd66998: data = 8'h05;
      17'd66999: data = 8'h01;
      17'd67000: data = 8'h02;
      17'd67001: data = 8'h01;
      17'd67002: data = 8'h01;
      17'd67003: data = 8'h0a;
      17'd67004: data = 8'h09;
      17'd67005: data = 8'h0c;
      17'd67006: data = 8'h0c;
      17'd67007: data = 8'h0a;
      17'd67008: data = 8'h0e;
      17'd67009: data = 8'h05;
      17'd67010: data = 8'h13;
      17'd67011: data = 8'h11;
      17'd67012: data = 8'h0a;
      17'd67013: data = 8'h11;
      17'd67014: data = 8'h0c;
      17'd67015: data = 8'h16;
      17'd67016: data = 8'h0c;
      17'd67017: data = 8'h12;
      17'd67018: data = 8'h12;
      17'd67019: data = 8'h0c;
      17'd67020: data = 8'h0e;
      17'd67021: data = 8'h09;
      17'd67022: data = 8'h0a;
      17'd67023: data = 8'h0c;
      17'd67024: data = 8'h0a;
      17'd67025: data = 8'h0d;
      17'd67026: data = 8'h13;
      17'd67027: data = 8'h0a;
      17'd67028: data = 8'h11;
      17'd67029: data = 8'h0d;
      17'd67030: data = 8'h05;
      17'd67031: data = 8'h06;
      17'd67032: data = 8'h09;
      17'd67033: data = 8'h0c;
      17'd67034: data = 8'h06;
      17'd67035: data = 8'h0d;
      17'd67036: data = 8'h09;
      17'd67037: data = 8'h09;
      17'd67038: data = 8'h0a;
      17'd67039: data = 8'h06;
      17'd67040: data = 8'h0a;
      17'd67041: data = 8'h09;
      17'd67042: data = 8'hfe;
      17'd67043: data = 8'hfd;
      17'd67044: data = 8'hfc;
      17'd67045: data = 8'hf9;
      17'd67046: data = 8'h02;
      17'd67047: data = 8'hfc;
      17'd67048: data = 8'h01;
      17'd67049: data = 8'h06;
      17'd67050: data = 8'h05;
      17'd67051: data = 8'h0e;
      17'd67052: data = 8'h1a;
      17'd67053: data = 8'h23;
      17'd67054: data = 8'h1f;
      17'd67055: data = 8'h1c;
      17'd67056: data = 8'h0a;
      17'd67057: data = 8'h02;
      17'd67058: data = 8'hfe;
      17'd67059: data = 8'hf9;
      17'd67060: data = 8'h02;
      17'd67061: data = 8'h0a;
      17'd67062: data = 8'h0a;
      17'd67063: data = 8'h11;
      17'd67064: data = 8'h12;
      17'd67065: data = 8'h06;
      17'd67066: data = 8'h19;
      17'd67067: data = 8'h1b;
      17'd67068: data = 8'h16;
      17'd67069: data = 8'h1a;
      17'd67070: data = 8'h11;
      17'd67071: data = 8'h0a;
      17'd67072: data = 8'h04;
      17'd67073: data = 8'h00;
      17'd67074: data = 8'h01;
      17'd67075: data = 8'h09;
      17'd67076: data = 8'h00;
      17'd67077: data = 8'hf9;
      17'd67078: data = 8'hf2;
      17'd67079: data = 8'he7;
      17'd67080: data = 8'hec;
      17'd67081: data = 8'hfa;
      17'd67082: data = 8'h02;
      17'd67083: data = 8'h05;
      17'd67084: data = 8'h09;
      17'd67085: data = 8'hfa;
      17'd67086: data = 8'hf1;
      17'd67087: data = 8'he9;
      17'd67088: data = 8'he3;
      17'd67089: data = 8'he9;
      17'd67090: data = 8'he2;
      17'd67091: data = 8'hda;
      17'd67092: data = 8'hd6;
      17'd67093: data = 8'hd6;
      17'd67094: data = 8'hd6;
      17'd67095: data = 8'he0;
      17'd67096: data = 8'he9;
      17'd67097: data = 8'hef;
      17'd67098: data = 8'hf1;
      17'd67099: data = 8'he9;
      17'd67100: data = 8'he5;
      17'd67101: data = 8'he5;
      17'd67102: data = 8'heb;
      17'd67103: data = 8'hec;
      17'd67104: data = 8'hf2;
      17'd67105: data = 8'hf2;
      17'd67106: data = 8'hf1;
      17'd67107: data = 8'heb;
      17'd67108: data = 8'he2;
      17'd67109: data = 8'he7;
      17'd67110: data = 8'hef;
      17'd67111: data = 8'hfa;
      17'd67112: data = 8'h01;
      17'd67113: data = 8'h05;
      17'd67114: data = 8'h0a;
      17'd67115: data = 8'h0e;
      17'd67116: data = 8'h12;
      17'd67117: data = 8'h11;
      17'd67118: data = 8'h19;
      17'd67119: data = 8'h13;
      17'd67120: data = 8'h11;
      17'd67121: data = 8'h0a;
      17'd67122: data = 8'h06;
      17'd67123: data = 8'h0a;
      17'd67124: data = 8'h0d;
      17'd67125: data = 8'h15;
      17'd67126: data = 8'h19;
      17'd67127: data = 8'h1c;
      17'd67128: data = 8'h19;
      17'd67129: data = 8'h1a;
      17'd67130: data = 8'h19;
      17'd67131: data = 8'h16;
      17'd67132: data = 8'h1a;
      17'd67133: data = 8'h16;
      17'd67134: data = 8'h19;
      17'd67135: data = 8'h15;
      17'd67136: data = 8'h11;
      17'd67137: data = 8'h0a;
      17'd67138: data = 8'h05;
      17'd67139: data = 8'hfd;
      17'd67140: data = 8'hfd;
      17'd67141: data = 8'hfc;
      17'd67142: data = 8'hf5;
      17'd67143: data = 8'hfa;
      17'd67144: data = 8'hfc;
      17'd67145: data = 8'hfe;
      17'd67146: data = 8'hfc;
      17'd67147: data = 8'hfc;
      17'd67148: data = 8'hf5;
      17'd67149: data = 8'hf1;
      17'd67150: data = 8'hed;
      17'd67151: data = 8'he4;
      17'd67152: data = 8'he4;
      17'd67153: data = 8'hde;
      17'd67154: data = 8'hdb;
      17'd67155: data = 8'hde;
      17'd67156: data = 8'hde;
      17'd67157: data = 8'he0;
      17'd67158: data = 8'he2;
      17'd67159: data = 8'hde;
      17'd67160: data = 8'hdc;
      17'd67161: data = 8'hde;
      17'd67162: data = 8'hdc;
      17'd67163: data = 8'hdc;
      17'd67164: data = 8'hde;
      17'd67165: data = 8'he0;
      17'd67166: data = 8'he0;
      17'd67167: data = 8'he4;
      17'd67168: data = 8'he3;
      17'd67169: data = 8'hdc;
      17'd67170: data = 8'he2;
      17'd67171: data = 8'he2;
      17'd67172: data = 8'he2;
      17'd67173: data = 8'he3;
      17'd67174: data = 8'he9;
      17'd67175: data = 8'hf1;
      17'd67176: data = 8'hef;
      17'd67177: data = 8'hf5;
      17'd67178: data = 8'hfc;
      17'd67179: data = 8'hfe;
      17'd67180: data = 8'hfe;
      17'd67181: data = 8'hfd;
      17'd67182: data = 8'hfd;
      17'd67183: data = 8'hfc;
      17'd67184: data = 8'hfc;
      17'd67185: data = 8'hfe;
      17'd67186: data = 8'h02;
      17'd67187: data = 8'h05;
      17'd67188: data = 8'h06;
      17'd67189: data = 8'h09;
      17'd67190: data = 8'h05;
      17'd67191: data = 8'h02;
      17'd67192: data = 8'h06;
      17'd67193: data = 8'h06;
      17'd67194: data = 8'h0a;
      17'd67195: data = 8'h0e;
      17'd67196: data = 8'h12;
      17'd67197: data = 8'h12;
      17'd67198: data = 8'h0c;
      17'd67199: data = 8'h0a;
      17'd67200: data = 8'h09;
      17'd67201: data = 8'h04;
      17'd67202: data = 8'h01;
      17'd67203: data = 8'h00;
      17'd67204: data = 8'hfd;
      17'd67205: data = 8'hfe;
      17'd67206: data = 8'hfe;
      17'd67207: data = 8'hfe;
      17'd67208: data = 8'h01;
      17'd67209: data = 8'h02;
      17'd67210: data = 8'h01;
      17'd67211: data = 8'h00;
      17'd67212: data = 8'hfd;
      17'd67213: data = 8'hf9;
      17'd67214: data = 8'hfc;
      17'd67215: data = 8'hfa;
      17'd67216: data = 8'hfc;
      17'd67217: data = 8'hfc;
      17'd67218: data = 8'hf6;
      17'd67219: data = 8'hf5;
      17'd67220: data = 8'hf2;
      17'd67221: data = 8'hf2;
      17'd67222: data = 8'hf4;
      17'd67223: data = 8'hf6;
      17'd67224: data = 8'hfa;
      17'd67225: data = 8'hfc;
      17'd67226: data = 8'hfc;
      17'd67227: data = 8'hfc;
      17'd67228: data = 8'hfd;
      17'd67229: data = 8'hfe;
      17'd67230: data = 8'hfd;
      17'd67231: data = 8'hfc;
      17'd67232: data = 8'hfc;
      17'd67233: data = 8'hfd;
      17'd67234: data = 8'hfe;
      17'd67235: data = 8'hfe;
      17'd67236: data = 8'h02;
      17'd67237: data = 8'h05;
      17'd67238: data = 8'h09;
      17'd67239: data = 8'h0a;
      17'd67240: data = 8'h0a;
      17'd67241: data = 8'h0c;
      17'd67242: data = 8'h0a;
      17'd67243: data = 8'h0d;
      17'd67244: data = 8'h11;
      17'd67245: data = 8'h0c;
      17'd67246: data = 8'h0e;
      17'd67247: data = 8'h0d;
      17'd67248: data = 8'h0e;
      17'd67249: data = 8'h0a;
      17'd67250: data = 8'h04;
      17'd67251: data = 8'h12;
      17'd67252: data = 8'h0c;
      17'd67253: data = 8'h13;
      17'd67254: data = 8'h13;
      17'd67255: data = 8'h13;
      17'd67256: data = 8'h15;
      17'd67257: data = 8'h13;
      17'd67258: data = 8'h19;
      17'd67259: data = 8'h0c;
      17'd67260: data = 8'h0d;
      17'd67261: data = 8'h04;
      17'd67262: data = 8'h06;
      17'd67263: data = 8'h02;
      17'd67264: data = 8'h06;
      17'd67265: data = 8'h04;
      17'd67266: data = 8'h15;
      17'd67267: data = 8'h05;
      17'd67268: data = 8'h05;
      17'd67269: data = 8'h12;
      17'd67270: data = 8'hfe;
      17'd67271: data = 8'h0d;
      17'd67272: data = 8'hfc;
      17'd67273: data = 8'h0c;
      17'd67274: data = 8'h01;
      17'd67275: data = 8'h02;
      17'd67276: data = 8'h05;
      17'd67277: data = 8'h01;
      17'd67278: data = 8'h05;
      17'd67279: data = 8'hfa;
      17'd67280: data = 8'hfc;
      17'd67281: data = 8'hfa;
      17'd67282: data = 8'hf9;
      17'd67283: data = 8'hf9;
      17'd67284: data = 8'h0a;
      17'd67285: data = 8'h02;
      17'd67286: data = 8'h13;
      17'd67287: data = 8'h0d;
      17'd67288: data = 8'h11;
      17'd67289: data = 8'h15;
      17'd67290: data = 8'h01;
      17'd67291: data = 8'h13;
      17'd67292: data = 8'h02;
      17'd67293: data = 8'h02;
      17'd67294: data = 8'h01;
      17'd67295: data = 8'h02;
      17'd67296: data = 8'h02;
      17'd67297: data = 8'h04;
      17'd67298: data = 8'h0d;
      17'd67299: data = 8'h11;
      17'd67300: data = 8'h1a;
      17'd67301: data = 8'h11;
      17'd67302: data = 8'h15;
      17'd67303: data = 8'h15;
      17'd67304: data = 8'h13;
      17'd67305: data = 8'h11;
      17'd67306: data = 8'h1c;
      17'd67307: data = 8'h12;
      17'd67308: data = 8'h13;
      17'd67309: data = 8'h11;
      17'd67310: data = 8'h06;
      17'd67311: data = 8'h09;
      17'd67312: data = 8'h00;
      17'd67313: data = 8'h0c;
      17'd67314: data = 8'h04;
      17'd67315: data = 8'h0a;
      17'd67316: data = 8'h02;
      17'd67317: data = 8'h01;
      17'd67318: data = 8'h01;
      17'd67319: data = 8'h01;
      17'd67320: data = 8'h09;
      17'd67321: data = 8'h0a;
      17'd67322: data = 8'h0c;
      17'd67323: data = 8'h05;
      17'd67324: data = 8'hfd;
      17'd67325: data = 8'hef;
      17'd67326: data = 8'hed;
      17'd67327: data = 8'he2;
      17'd67328: data = 8'heb;
      17'd67329: data = 8'he7;
      17'd67330: data = 8'hed;
      17'd67331: data = 8'heb;
      17'd67332: data = 8'he2;
      17'd67333: data = 8'he7;
      17'd67334: data = 8'hde;
      17'd67335: data = 8'heb;
      17'd67336: data = 8'heb;
      17'd67337: data = 8'hf1;
      17'd67338: data = 8'hec;
      17'd67339: data = 8'he3;
      17'd67340: data = 8'he2;
      17'd67341: data = 8'hd8;
      17'd67342: data = 8'hdb;
      17'd67343: data = 8'he2;
      17'd67344: data = 8'he4;
      17'd67345: data = 8'he2;
      17'd67346: data = 8'hde;
      17'd67347: data = 8'hd3;
      17'd67348: data = 8'hd8;
      17'd67349: data = 8'hdb;
      17'd67350: data = 8'he9;
      17'd67351: data = 8'hf5;
      17'd67352: data = 8'hfa;
      17'd67353: data = 8'hfc;
      17'd67354: data = 8'hf2;
      17'd67355: data = 8'hf5;
      17'd67356: data = 8'hf1;
      17'd67357: data = 8'hfc;
      17'd67358: data = 8'h01;
      17'd67359: data = 8'h04;
      17'd67360: data = 8'h05;
      17'd67361: data = 8'hfe;
      17'd67362: data = 8'h04;
      17'd67363: data = 8'h00;
      17'd67364: data = 8'h06;
      17'd67365: data = 8'h12;
      17'd67366: data = 8'h15;
      17'd67367: data = 8'h1a;
      17'd67368: data = 8'h16;
      17'd67369: data = 8'h15;
      17'd67370: data = 8'h19;
      17'd67371: data = 8'h1b;
      17'd67372: data = 8'h23;
      17'd67373: data = 8'h26;
      17'd67374: data = 8'h24;
      17'd67375: data = 8'h1c;
      17'd67376: data = 8'h11;
      17'd67377: data = 8'h0e;
      17'd67378: data = 8'h06;
      17'd67379: data = 8'h0e;
      17'd67380: data = 8'h13;
      17'd67381: data = 8'h13;
      17'd67382: data = 8'h15;
      17'd67383: data = 8'h0e;
      17'd67384: data = 8'h0d;
      17'd67385: data = 8'h0a;
      17'd67386: data = 8'h09;
      17'd67387: data = 8'h0a;
      17'd67388: data = 8'h05;
      17'd67389: data = 8'h02;
      17'd67390: data = 8'hfd;
      17'd67391: data = 8'hf5;
      17'd67392: data = 8'hef;
      17'd67393: data = 8'hec;
      17'd67394: data = 8'hec;
      17'd67395: data = 8'hec;
      17'd67396: data = 8'he9;
      17'd67397: data = 8'he4;
      17'd67398: data = 8'hdc;
      17'd67399: data = 8'hdc;
      17'd67400: data = 8'hdc;
      17'd67401: data = 8'he0;
      17'd67402: data = 8'he4;
      17'd67403: data = 8'he5;
      17'd67404: data = 8'he7;
      17'd67405: data = 8'he5;
      17'd67406: data = 8'he2;
      17'd67407: data = 8'hdb;
      17'd67408: data = 8'hd6;
      17'd67409: data = 8'hd6;
      17'd67410: data = 8'hd8;
      17'd67411: data = 8'hd8;
      17'd67412: data = 8'hd8;
      17'd67413: data = 8'hdb;
      17'd67414: data = 8'he0;
      17'd67415: data = 8'he4;
      17'd67416: data = 8'heb;
      17'd67417: data = 8'hef;
      17'd67418: data = 8'hf1;
      17'd67419: data = 8'hf1;
      17'd67420: data = 8'hef;
      17'd67421: data = 8'hf1;
      17'd67422: data = 8'hf2;
      17'd67423: data = 8'hf9;
      17'd67424: data = 8'hfc;
      17'd67425: data = 8'hfd;
      17'd67426: data = 8'hfe;
      17'd67427: data = 8'hfc;
      17'd67428: data = 8'hfc;
      17'd67429: data = 8'hf9;
      17'd67430: data = 8'hfc;
      17'd67431: data = 8'h02;
      17'd67432: data = 8'h0a;
      17'd67433: data = 8'h0d;
      17'd67434: data = 8'h15;
      17'd67435: data = 8'h19;
      17'd67436: data = 8'h19;
      17'd67437: data = 8'h19;
      17'd67438: data = 8'h13;
      17'd67439: data = 8'h12;
      17'd67440: data = 8'h0e;
      17'd67441: data = 8'h0a;
      17'd67442: data = 8'h09;
      17'd67443: data = 8'h09;
      17'd67444: data = 8'h05;
      17'd67445: data = 8'h06;
      17'd67446: data = 8'h06;
      17'd67447: data = 8'h06;
      17'd67448: data = 8'h09;
      17'd67449: data = 8'h04;
      17'd67450: data = 8'h05;
      17'd67451: data = 8'h04;
      17'd67452: data = 8'h01;
      17'd67453: data = 8'h02;
      17'd67454: data = 8'h02;
      17'd67455: data = 8'h01;
      17'd67456: data = 8'hfd;
      17'd67457: data = 8'hf9;
      17'd67458: data = 8'hf1;
      17'd67459: data = 8'heb;
      17'd67460: data = 8'he5;
      17'd67461: data = 8'he5;
      17'd67462: data = 8'heb;
      17'd67463: data = 8'hed;
      17'd67464: data = 8'hf1;
      17'd67465: data = 8'hf4;
      17'd67466: data = 8'hf5;
      17'd67467: data = 8'hf5;
      17'd67468: data = 8'hf9;
      17'd67469: data = 8'hf5;
      17'd67470: data = 8'hf4;
      17'd67471: data = 8'hf2;
      17'd67472: data = 8'hef;
      17'd67473: data = 8'hf4;
      17'd67474: data = 8'hf4;
      17'd67475: data = 8'hf4;
      17'd67476: data = 8'hfa;
      17'd67477: data = 8'hfc;
      17'd67478: data = 8'hf9;
      17'd67479: data = 8'hfc;
      17'd67480: data = 8'hfa;
      17'd67481: data = 8'hfe;
      17'd67482: data = 8'h05;
      17'd67483: data = 8'h09;
      17'd67484: data = 8'h13;
      17'd67485: data = 8'h15;
      17'd67486: data = 8'h16;
      17'd67487: data = 8'h1a;
      17'd67488: data = 8'h11;
      17'd67489: data = 8'h13;
      17'd67490: data = 8'h12;
      17'd67491: data = 8'h09;
      17'd67492: data = 8'h15;
      17'd67493: data = 8'h12;
      17'd67494: data = 8'h13;
      17'd67495: data = 8'h1c;
      17'd67496: data = 8'h1a;
      17'd67497: data = 8'h1b;
      17'd67498: data = 8'h1f;
      17'd67499: data = 8'h1c;
      17'd67500: data = 8'h1b;
      17'd67501: data = 8'h1e;
      17'd67502: data = 8'h13;
      17'd67503: data = 8'h19;
      17'd67504: data = 8'h1a;
      17'd67505: data = 8'h16;
      17'd67506: data = 8'h16;
      17'd67507: data = 8'h1b;
      17'd67508: data = 8'h0e;
      17'd67509: data = 8'h0e;
      17'd67510: data = 8'h0a;
      17'd67511: data = 8'h01;
      17'd67512: data = 8'h06;
      17'd67513: data = 8'h04;
      17'd67514: data = 8'h04;
      17'd67515: data = 8'h0c;
      17'd67516: data = 8'h0a;
      17'd67517: data = 8'h05;
      17'd67518: data = 8'h0a;
      17'd67519: data = 8'h00;
      17'd67520: data = 8'h04;
      17'd67521: data = 8'hfe;
      17'd67522: data = 8'hfd;
      17'd67523: data = 8'hfe;
      17'd67524: data = 8'h02;
      17'd67525: data = 8'h02;
      17'd67526: data = 8'h02;
      17'd67527: data = 8'h04;
      17'd67528: data = 8'h09;
      17'd67529: data = 8'h01;
      17'd67530: data = 8'hfe;
      17'd67531: data = 8'h06;
      17'd67532: data = 8'hfe;
      17'd67533: data = 8'h05;
      17'd67534: data = 8'h06;
      17'd67535: data = 8'h0a;
      17'd67536: data = 8'h11;
      17'd67537: data = 8'h0d;
      17'd67538: data = 8'h13;
      17'd67539: data = 8'h1a;
      17'd67540: data = 8'h15;
      17'd67541: data = 8'h0c;
      17'd67542: data = 8'h06;
      17'd67543: data = 8'hfc;
      17'd67544: data = 8'hf4;
      17'd67545: data = 8'hfd;
      17'd67546: data = 8'h05;
      17'd67547: data = 8'h19;
      17'd67548: data = 8'h2c;
      17'd67549: data = 8'h2f;
      17'd67550: data = 8'h2f;
      17'd67551: data = 8'h27;
      17'd67552: data = 8'h13;
      17'd67553: data = 8'h16;
      17'd67554: data = 8'h13;
      17'd67555: data = 8'h12;
      17'd67556: data = 8'h1b;
      17'd67557: data = 8'h12;
      17'd67558: data = 8'h06;
      17'd67559: data = 8'h04;
      17'd67560: data = 8'hfe;
      17'd67561: data = 8'h01;
      17'd67562: data = 8'h0e;
      17'd67563: data = 8'h06;
      17'd67564: data = 8'h09;
      17'd67565: data = 8'h09;
      17'd67566: data = 8'hfd;
      17'd67567: data = 8'h05;
      17'd67568: data = 8'h0a;
      17'd67569: data = 8'h0e;
      17'd67570: data = 8'h16;
      17'd67571: data = 8'h06;
      17'd67572: data = 8'hf6;
      17'd67573: data = 8'he3;
      17'd67574: data = 8'hd2;
      17'd67575: data = 8'hd1;
      17'd67576: data = 8'hd6;
      17'd67577: data = 8'he4;
      17'd67578: data = 8'hec;
      17'd67579: data = 8'hf5;
      17'd67580: data = 8'hef;
      17'd67581: data = 8'he7;
      17'd67582: data = 8'he3;
      17'd67583: data = 8'hdc;
      17'd67584: data = 8'he5;
      17'd67585: data = 8'he5;
      17'd67586: data = 8'he2;
      17'd67587: data = 8'he4;
      17'd67588: data = 8'hda;
      17'd67589: data = 8'hd8;
      17'd67590: data = 8'hd8;
      17'd67591: data = 8'hd5;
      17'd67592: data = 8'hdb;
      17'd67593: data = 8'hda;
      17'd67594: data = 8'hd6;
      17'd67595: data = 8'hdb;
      17'd67596: data = 8'he0;
      17'd67597: data = 8'he9;
      17'd67598: data = 8'hf5;
      17'd67599: data = 8'h02;
      17'd67600: data = 8'h09;
      17'd67601: data = 8'h0c;
      17'd67602: data = 8'h04;
      17'd67603: data = 8'hfa;
      17'd67604: data = 8'hf4;
      17'd67605: data = 8'hf1;
      17'd67606: data = 8'hf5;
      17'd67607: data = 8'hfd;
      17'd67608: data = 8'h04;
      17'd67609: data = 8'h0d;
      17'd67610: data = 8'h15;
      17'd67611: data = 8'h13;
      17'd67612: data = 8'h15;
      17'd67613: data = 8'h16;
      17'd67614: data = 8'h19;
      17'd67615: data = 8'h1a;
      17'd67616: data = 8'h1c;
      17'd67617: data = 8'h1e;
      17'd67618: data = 8'h24;
      17'd67619: data = 8'h22;
      17'd67620: data = 8'h22;
      17'd67621: data = 8'h1e;
      17'd67622: data = 8'h15;
      17'd67623: data = 8'h0e;
      17'd67624: data = 8'h09;
      17'd67625: data = 8'h06;
      17'd67626: data = 8'h0a;
      17'd67627: data = 8'h0d;
      17'd67628: data = 8'h15;
      17'd67629: data = 8'h16;
      17'd67630: data = 8'h19;
      17'd67631: data = 8'h19;
      17'd67632: data = 8'h15;
      17'd67633: data = 8'h0e;
      17'd67634: data = 8'h04;
      17'd67635: data = 8'hfd;
      17'd67636: data = 8'hf2;
      17'd67637: data = 8'hed;
      17'd67638: data = 8'heb;
      17'd67639: data = 8'heb;
      17'd67640: data = 8'hf1;
      17'd67641: data = 8'hf1;
      17'd67642: data = 8'heb;
      17'd67643: data = 8'he5;
      17'd67644: data = 8'he0;
      17'd67645: data = 8'he0;
      17'd67646: data = 8'he2;
      17'd67647: data = 8'he4;
      17'd67648: data = 8'he9;
      17'd67649: data = 8'hec;
      17'd67650: data = 8'he7;
      17'd67651: data = 8'he0;
      17'd67652: data = 8'hdc;
      17'd67653: data = 8'hd6;
      17'd67654: data = 8'hd3;
      17'd67655: data = 8'hd3;
      17'd67656: data = 8'hd3;
      17'd67657: data = 8'hd6;
      17'd67658: data = 8'hdc;
      17'd67659: data = 8'he0;
      17'd67660: data = 8'he9;
      17'd67661: data = 8'hf4;
      17'd67662: data = 8'hf6;
      17'd67663: data = 8'hf9;
      17'd67664: data = 8'hf5;
      17'd67665: data = 8'hed;
      17'd67666: data = 8'he9;
      17'd67667: data = 8'he5;
      17'd67668: data = 8'heb;
      17'd67669: data = 8'hf1;
      17'd67670: data = 8'hf5;
      17'd67671: data = 8'hfc;
      17'd67672: data = 8'h00;
      17'd67673: data = 8'h01;
      17'd67674: data = 8'h00;
      17'd67675: data = 8'h00;
      17'd67676: data = 8'h02;
      17'd67677: data = 8'h06;
      17'd67678: data = 8'h0c;
      17'd67679: data = 8'h12;
      17'd67680: data = 8'h15;
      17'd67681: data = 8'h13;
      17'd67682: data = 8'h13;
      17'd67683: data = 8'h0c;
      17'd67684: data = 8'h04;
      17'd67685: data = 8'h01;
      17'd67686: data = 8'hfd;
      17'd67687: data = 8'hfe;
      17'd67688: data = 8'h04;
      17'd67689: data = 8'h09;
      17'd67690: data = 8'h0d;
      17'd67691: data = 8'h12;
      17'd67692: data = 8'h12;
      17'd67693: data = 8'h12;
      17'd67694: data = 8'h0d;
      17'd67695: data = 8'h06;
      17'd67696: data = 8'h02;
      17'd67697: data = 8'hfd;
      17'd67698: data = 8'hf9;
      17'd67699: data = 8'hf9;
      17'd67700: data = 8'hf6;
      17'd67701: data = 8'hf6;
      17'd67702: data = 8'hfa;
      17'd67703: data = 8'hf5;
      17'd67704: data = 8'hf2;
      17'd67705: data = 8'hef;
      17'd67706: data = 8'heb;
      17'd67707: data = 8'hec;
      17'd67708: data = 8'hef;
      17'd67709: data = 8'hf2;
      17'd67710: data = 8'hf9;
      17'd67711: data = 8'hfa;
      17'd67712: data = 8'hf9;
      17'd67713: data = 8'hf1;
      17'd67714: data = 8'he9;
      17'd67715: data = 8'he2;
      17'd67716: data = 8'he0;
      17'd67717: data = 8'hde;
      17'd67718: data = 8'he3;
      17'd67719: data = 8'hec;
      17'd67720: data = 8'hf1;
      17'd67721: data = 8'hf6;
      17'd67722: data = 8'hfa;
      17'd67723: data = 8'hfc;
      17'd67724: data = 8'hfc;
      17'd67725: data = 8'hfa;
      17'd67726: data = 8'hfc;
      17'd67727: data = 8'hfa;
      17'd67728: data = 8'hfa;
      17'd67729: data = 8'hfc;
      17'd67730: data = 8'h00;
      17'd67731: data = 8'h04;
      17'd67732: data = 8'h0a;
      17'd67733: data = 8'h0a;
      17'd67734: data = 8'h09;
      17'd67735: data = 8'h09;
      17'd67736: data = 8'h05;
      17'd67737: data = 8'h09;
      17'd67738: data = 8'h0e;
      17'd67739: data = 8'h13;
      17'd67740: data = 8'h1b;
      17'd67741: data = 8'h22;
      17'd67742: data = 8'h1e;
      17'd67743: data = 8'h1f;
      17'd67744: data = 8'h19;
      17'd67745: data = 8'h15;
      17'd67746: data = 8'h13;
      17'd67747: data = 8'h0e;
      17'd67748: data = 8'h11;
      17'd67749: data = 8'h0e;
      17'd67750: data = 8'h12;
      17'd67751: data = 8'h16;
      17'd67752: data = 8'h1c;
      17'd67753: data = 8'h19;
      17'd67754: data = 8'h13;
      17'd67755: data = 8'h13;
      17'd67756: data = 8'h11;
      17'd67757: data = 8'h15;
      17'd67758: data = 8'h0d;
      17'd67759: data = 8'h12;
      17'd67760: data = 8'h0d;
      17'd67761: data = 8'h0c;
      17'd67762: data = 8'h0e;
      17'd67763: data = 8'h0a;
      17'd67764: data = 8'hfd;
      17'd67765: data = 8'hfd;
      17'd67766: data = 8'hfc;
      17'd67767: data = 8'hfa;
      17'd67768: data = 8'h01;
      17'd67769: data = 8'h06;
      17'd67770: data = 8'h09;
      17'd67771: data = 8'hfe;
      17'd67772: data = 8'hfe;
      17'd67773: data = 8'h06;
      17'd67774: data = 8'h05;
      17'd67775: data = 8'h09;
      17'd67776: data = 8'h0e;
      17'd67777: data = 8'h0c;
      17'd67778: data = 8'h02;
      17'd67779: data = 8'h01;
      17'd67780: data = 8'h02;
      17'd67781: data = 8'h00;
      17'd67782: data = 8'h04;
      17'd67783: data = 8'h0a;
      17'd67784: data = 8'h09;
      17'd67785: data = 8'h15;
      17'd67786: data = 8'h19;
      17'd67787: data = 8'h0a;
      17'd67788: data = 8'h0e;
      17'd67789: data = 8'h0c;
      17'd67790: data = 8'h0e;
      17'd67791: data = 8'h11;
      17'd67792: data = 8'h11;
      17'd67793: data = 8'h12;
      17'd67794: data = 8'h16;
      17'd67795: data = 8'h0e;
      17'd67796: data = 8'h0d;
      17'd67797: data = 8'h0e;
      17'd67798: data = 8'h0a;
      17'd67799: data = 8'h02;
      17'd67800: data = 8'h02;
      17'd67801: data = 8'h05;
      17'd67802: data = 8'h06;
      17'd67803: data = 8'h0c;
      17'd67804: data = 8'h0d;
      17'd67805: data = 8'h11;
      17'd67806: data = 8'h0d;
      17'd67807: data = 8'h0c;
      17'd67808: data = 8'h06;
      17'd67809: data = 8'h04;
      17'd67810: data = 8'hfe;
      17'd67811: data = 8'hfd;
      17'd67812: data = 8'hf6;
      17'd67813: data = 8'hf5;
      17'd67814: data = 8'hf5;
      17'd67815: data = 8'hf4;
      17'd67816: data = 8'hf4;
      17'd67817: data = 8'hf2;
      17'd67818: data = 8'hf4;
      17'd67819: data = 8'hf6;
      17'd67820: data = 8'hf6;
      17'd67821: data = 8'hf6;
      17'd67822: data = 8'hf9;
      17'd67823: data = 8'hf6;
      17'd67824: data = 8'hf5;
      17'd67825: data = 8'hf4;
      17'd67826: data = 8'hf1;
      17'd67827: data = 8'hef;
      17'd67828: data = 8'hec;
      17'd67829: data = 8'hed;
      17'd67830: data = 8'hed;
      17'd67831: data = 8'hec;
      17'd67832: data = 8'hed;
      17'd67833: data = 8'hed;
      17'd67834: data = 8'hed;
      17'd67835: data = 8'hf1;
      17'd67836: data = 8'hf5;
      17'd67837: data = 8'hf5;
      17'd67838: data = 8'hfa;
      17'd67839: data = 8'hfa;
      17'd67840: data = 8'hf5;
      17'd67841: data = 8'hf6;
      17'd67842: data = 8'hf5;
      17'd67843: data = 8'hf2;
      17'd67844: data = 8'hf1;
      17'd67845: data = 8'hef;
      17'd67846: data = 8'hef;
      17'd67847: data = 8'hed;
      17'd67848: data = 8'hef;
      17'd67849: data = 8'hef;
      17'd67850: data = 8'hf1;
      17'd67851: data = 8'hf2;
      17'd67852: data = 8'hf4;
      17'd67853: data = 8'hfc;
      17'd67854: data = 8'hfe;
      17'd67855: data = 8'h00;
      17'd67856: data = 8'h02;
      17'd67857: data = 8'h00;
      17'd67858: data = 8'h00;
      17'd67859: data = 8'hfc;
      17'd67860: data = 8'hf9;
      17'd67861: data = 8'hf9;
      17'd67862: data = 8'hf6;
      17'd67863: data = 8'hfa;
      17'd67864: data = 8'hf9;
      17'd67865: data = 8'hfd;
      17'd67866: data = 8'h00;
      17'd67867: data = 8'h04;
      17'd67868: data = 8'h05;
      17'd67869: data = 8'h05;
      17'd67870: data = 8'h04;
      17'd67871: data = 8'h04;
      17'd67872: data = 8'h05;
      17'd67873: data = 8'h04;
      17'd67874: data = 8'h04;
      17'd67875: data = 8'h01;
      17'd67876: data = 8'h01;
      17'd67877: data = 8'h01;
      17'd67878: data = 8'hfe;
      17'd67879: data = 8'hfe;
      17'd67880: data = 8'hfe;
      17'd67881: data = 8'hfe;
      17'd67882: data = 8'h00;
      17'd67883: data = 8'h01;
      17'd67884: data = 8'h01;
      17'd67885: data = 8'h01;
      17'd67886: data = 8'h00;
      17'd67887: data = 8'hfe;
      17'd67888: data = 8'hfe;
      17'd67889: data = 8'hfd;
      17'd67890: data = 8'hfd;
      17'd67891: data = 8'hfd;
      17'd67892: data = 8'hfa;
      17'd67893: data = 8'hf6;
      17'd67894: data = 8'hf5;
      17'd67895: data = 8'hf6;
      17'd67896: data = 8'hf9;
      17'd67897: data = 8'hf9;
      17'd67898: data = 8'hfa;
      17'd67899: data = 8'hfc;
      17'd67900: data = 8'hfe;
      17'd67901: data = 8'hfd;
      17'd67902: data = 8'hfc;
      17'd67903: data = 8'hfd;
      17'd67904: data = 8'hfc;
      17'd67905: data = 8'hfa;
      17'd67906: data = 8'hf6;
      17'd67907: data = 8'hf4;
      17'd67908: data = 8'hf4;
      17'd67909: data = 8'hf5;
      17'd67910: data = 8'hf9;
      17'd67911: data = 8'hfa;
      17'd67912: data = 8'hfe;
      17'd67913: data = 8'h00;
      17'd67914: data = 8'h00;
      17'd67915: data = 8'h01;
      17'd67916: data = 8'hfe;
      17'd67917: data = 8'hfe;
      17'd67918: data = 8'hfd;
      17'd67919: data = 8'hfc;
      17'd67920: data = 8'hfc;
      17'd67921: data = 8'hfa;
      17'd67922: data = 8'hfc;
      17'd67923: data = 8'hfd;
      17'd67924: data = 8'h01;
      17'd67925: data = 8'h00;
      17'd67926: data = 8'h00;
      17'd67927: data = 8'hfe;
      17'd67928: data = 8'hfd;
      17'd67929: data = 8'hfc;
      17'd67930: data = 8'hf9;
      17'd67931: data = 8'hf9;
      17'd67932: data = 8'hf9;
      17'd67933: data = 8'hf9;
      17'd67934: data = 8'hf9;
      17'd67935: data = 8'hfa;
      17'd67936: data = 8'hf9;
      17'd67937: data = 8'hfa;
      17'd67938: data = 8'hfd;
      17'd67939: data = 8'hfa;
      17'd67940: data = 8'hfa;
      17'd67941: data = 8'hf6;
      17'd67942: data = 8'hf5;
      17'd67943: data = 8'hf4;
      17'd67944: data = 8'hf2;
      17'd67945: data = 8'hf2;
      17'd67946: data = 8'hf4;
      17'd67947: data = 8'hf9;
      17'd67948: data = 8'hfa;
      17'd67949: data = 8'hfa;
      17'd67950: data = 8'hfa;
      17'd67951: data = 8'hfa;
      17'd67952: data = 8'hf6;
      17'd67953: data = 8'hf5;
      17'd67954: data = 8'hf6;
      17'd67955: data = 8'hf9;
      17'd67956: data = 8'hfa;
      17'd67957: data = 8'hfc;
      17'd67958: data = 8'hfc;
      17'd67959: data = 8'hfa;
      17'd67960: data = 8'hfd;
      17'd67961: data = 8'hfe;
      17'd67962: data = 8'hfe;
      17'd67963: data = 8'h00;
      17'd67964: data = 8'h00;
      17'd67965: data = 8'h00;
      17'd67966: data = 8'h00;
      17'd67967: data = 8'h01;
      17'd67968: data = 8'h02;
      17'd67969: data = 8'h02;
      17'd67970: data = 8'h05;
      17'd67971: data = 8'h05;
      17'd67972: data = 8'h05;
      17'd67973: data = 8'h09;
      17'd67974: data = 8'h05;
      17'd67975: data = 8'h09;
      17'd67976: data = 8'h06;
      17'd67977: data = 8'h05;
      17'd67978: data = 8'h06;
      17'd67979: data = 8'h05;
      17'd67980: data = 8'h06;
      17'd67981: data = 8'h06;
      17'd67982: data = 8'h09;
      17'd67983: data = 8'h09;
      17'd67984: data = 8'h0a;
      17'd67985: data = 8'h0c;
      17'd67986: data = 8'h0a;
      17'd67987: data = 8'h0a;
      17'd67988: data = 8'h0a;
      17'd67989: data = 8'h05;
      17'd67990: data = 8'h06;
      17'd67991: data = 8'h05;
      17'd67992: data = 8'h05;
      17'd67993: data = 8'h06;
      17'd67994: data = 8'h05;
      17'd67995: data = 8'h06;
      17'd67996: data = 8'h09;
      17'd67997: data = 8'h09;
      17'd67998: data = 8'h0a;
      17'd67999: data = 8'h0a;
      17'd68000: data = 8'h06;
      17'd68001: data = 8'h05;
      17'd68002: data = 8'h04;
      17'd68003: data = 8'h02;
      17'd68004: data = 8'h02;
      17'd68005: data = 8'h02;
      17'd68006: data = 8'h05;
      17'd68007: data = 8'h05;
      17'd68008: data = 8'h05;
      17'd68009: data = 8'h05;
      17'd68010: data = 8'h05;
      17'd68011: data = 8'h06;
      17'd68012: data = 8'h05;
      17'd68013: data = 8'h06;
      17'd68014: data = 8'h06;
      17'd68015: data = 8'h06;
      17'd68016: data = 8'h06;
      17'd68017: data = 8'h06;
      17'd68018: data = 8'h05;
      17'd68019: data = 8'h05;
      17'd68020: data = 8'h09;
      17'd68021: data = 8'h09;
      17'd68022: data = 8'h09;
      17'd68023: data = 8'h06;
      17'd68024: data = 8'h09;
      17'd68025: data = 8'h0a;
      17'd68026: data = 8'h0a;
      17'd68027: data = 8'h0c;
      17'd68028: data = 8'h0d;
      17'd68029: data = 8'h0e;
      17'd68030: data = 8'h11;
      17'd68031: data = 8'h0e;
      17'd68032: data = 8'h0d;
      17'd68033: data = 8'h0e;
      17'd68034: data = 8'h0d;
      17'd68035: data = 8'h0a;
      17'd68036: data = 8'h09;
      17'd68037: data = 8'h0a;
      17'd68038: data = 8'h0c;
      17'd68039: data = 8'h0a;
      17'd68040: data = 8'h0d;
      17'd68041: data = 8'h0d;
      17'd68042: data = 8'h0e;
      17'd68043: data = 8'h11;
      17'd68044: data = 8'h0e;
      17'd68045: data = 8'h11;
      17'd68046: data = 8'h0d;
      17'd68047: data = 8'h0a;
      17'd68048: data = 8'h0a;
      17'd68049: data = 8'h0a;
      17'd68050: data = 8'h09;
      17'd68051: data = 8'h06;
      17'd68052: data = 8'h06;
      17'd68053: data = 8'h06;
      17'd68054: data = 8'h05;
      17'd68055: data = 8'h05;
      17'd68056: data = 8'h06;
      17'd68057: data = 8'h05;
      17'd68058: data = 8'h06;
      17'd68059: data = 8'h05;
      17'd68060: data = 8'h04;
      17'd68061: data = 8'h05;
      17'd68062: data = 8'h02;
      17'd68063: data = 8'h01;
      17'd68064: data = 8'h01;
      17'd68065: data = 8'h00;
      17'd68066: data = 8'hfe;
      17'd68067: data = 8'hfd;
      17'd68068: data = 8'hfc;
      17'd68069: data = 8'hfc;
      17'd68070: data = 8'hfc;
      17'd68071: data = 8'hfc;
      17'd68072: data = 8'hfa;
      17'd68073: data = 8'hfa;
      17'd68074: data = 8'hf9;
      17'd68075: data = 8'hfa;
      17'd68076: data = 8'hfa;
      17'd68077: data = 8'hf9;
      17'd68078: data = 8'hf6;
      17'd68079: data = 8'hf5;
      17'd68080: data = 8'hf5;
      17'd68081: data = 8'hf5;
      17'd68082: data = 8'hf4;
      17'd68083: data = 8'hf1;
      17'd68084: data = 8'hf1;
      17'd68085: data = 8'hf4;
      17'd68086: data = 8'hf4;
      17'd68087: data = 8'hf5;
      17'd68088: data = 8'hf5;
      17'd68089: data = 8'hf6;
      17'd68090: data = 8'hf6;
      17'd68091: data = 8'hf5;
      17'd68092: data = 8'hf6;
      17'd68093: data = 8'hf5;
      17'd68094: data = 8'hf5;
      17'd68095: data = 8'hf6;
      17'd68096: data = 8'hf4;
      17'd68097: data = 8'hf2;
      17'd68098: data = 8'hf5;
      17'd68099: data = 8'hf5;
      17'd68100: data = 8'hf9;
      17'd68101: data = 8'hfa;
      17'd68102: data = 8'hfc;
      17'd68103: data = 8'hfa;
      17'd68104: data = 8'hf6;
      17'd68105: data = 8'hf6;
      17'd68106: data = 8'hf6;
      17'd68107: data = 8'hf6;
      17'd68108: data = 8'hf6;
      17'd68109: data = 8'hf9;
      17'd68110: data = 8'hf9;
      17'd68111: data = 8'hf6;
      17'd68112: data = 8'hf6;
      17'd68113: data = 8'hf6;
      17'd68114: data = 8'hf2;
      17'd68115: data = 8'hf4;
      17'd68116: data = 8'hf5;
      17'd68117: data = 8'hf5;
      17'd68118: data = 8'hf9;
      17'd68119: data = 8'hf9;
      17'd68120: data = 8'hf9;
      17'd68121: data = 8'hf6;
      17'd68122: data = 8'hf9;
      17'd68123: data = 8'hf5;
      17'd68124: data = 8'hf5;
      17'd68125: data = 8'hf5;
      17'd68126: data = 8'hf5;
      17'd68127: data = 8'hf5;
      17'd68128: data = 8'hf4;
      17'd68129: data = 8'hf4;
      17'd68130: data = 8'hf4;
      17'd68131: data = 8'hf6;
      17'd68132: data = 8'hf6;
      17'd68133: data = 8'hf4;
      17'd68134: data = 8'hf5;
      17'd68135: data = 8'hf6;
      17'd68136: data = 8'hf6;
      17'd68137: data = 8'hf5;
      17'd68138: data = 8'hf6;
      17'd68139: data = 8'hf6;
      17'd68140: data = 8'hf6;
      17'd68141: data = 8'hf6;
      17'd68142: data = 8'hf4;
      17'd68143: data = 8'hf4;
      17'd68144: data = 8'hf4;
      17'd68145: data = 8'hf4;
      17'd68146: data = 8'hf5;
      17'd68147: data = 8'hf6;
      17'd68148: data = 8'hf6;
      17'd68149: data = 8'hf9;
      17'd68150: data = 8'hf6;
      17'd68151: data = 8'hfa;
      17'd68152: data = 8'hfc;
      17'd68153: data = 8'hf9;
      17'd68154: data = 8'hf9;
      17'd68155: data = 8'hfa;
      17'd68156: data = 8'hfa;
      17'd68157: data = 8'hf9;
      17'd68158: data = 8'hfc;
      17'd68159: data = 8'hfc;
      17'd68160: data = 8'hfd;
      17'd68161: data = 8'hfe;
      17'd68162: data = 8'h01;
      17'd68163: data = 8'h01;
      17'd68164: data = 8'h00;
      17'd68165: data = 8'h00;
      17'd68166: data = 8'hfe;
      17'd68167: data = 8'h00;
      17'd68168: data = 8'h01;
      17'd68169: data = 8'h01;
      17'd68170: data = 8'h02;
      17'd68171: data = 8'h05;
      17'd68172: data = 8'h04;
      17'd68173: data = 8'h01;
      17'd68174: data = 8'h02;
      17'd68175: data = 8'h01;
      17'd68176: data = 8'h01;
      17'd68177: data = 8'h02;
      17'd68178: data = 8'h04;
      17'd68179: data = 8'h05;
      17'd68180: data = 8'h04;
      17'd68181: data = 8'h04;
      17'd68182: data = 8'h04;
      17'd68183: data = 8'h05;
      17'd68184: data = 8'h05;
      17'd68185: data = 8'h04;
      17'd68186: data = 8'h01;
      17'd68187: data = 8'h04;
      17'd68188: data = 8'h02;
      17'd68189: data = 8'h02;
      17'd68190: data = 8'h02;
      17'd68191: data = 8'h02;
      17'd68192: data = 8'h01;
      17'd68193: data = 8'h00;
      17'd68194: data = 8'h01;
      17'd68195: data = 8'h01;
      17'd68196: data = 8'h01;
      17'd68197: data = 8'h01;
      17'd68198: data = 8'h02;
      17'd68199: data = 8'h02;
      17'd68200: data = 8'h00;
      17'd68201: data = 8'h01;
      17'd68202: data = 8'h00;
      17'd68203: data = 8'h00;
      17'd68204: data = 8'h01;
      17'd68205: data = 8'h00;
      17'd68206: data = 8'h01;
      17'd68207: data = 8'h01;
      17'd68208: data = 8'h00;
      17'd68209: data = 8'h01;
      17'd68210: data = 8'h02;
      17'd68211: data = 8'h04;
      17'd68212: data = 8'h04;
      17'd68213: data = 8'h04;
      17'd68214: data = 8'h05;
      17'd68215: data = 8'h02;
      17'd68216: data = 8'h02;
      17'd68217: data = 8'h01;
      17'd68218: data = 8'h02;
      17'd68219: data = 8'h04;
      17'd68220: data = 8'h04;
      17'd68221: data = 8'h04;
      17'd68222: data = 8'h04;
      17'd68223: data = 8'h06;
      17'd68224: data = 8'h04;
      17'd68225: data = 8'h04;
      17'd68226: data = 8'h04;
      17'd68227: data = 8'h04;
      17'd68228: data = 8'h04;
      17'd68229: data = 8'h02;
      17'd68230: data = 8'h05;
      17'd68231: data = 8'h05;
      17'd68232: data = 8'h02;
      17'd68233: data = 8'h04;
      17'd68234: data = 8'h04;
      17'd68235: data = 8'h01;
      17'd68236: data = 8'h02;
      17'd68237: data = 8'h04;
      17'd68238: data = 8'h02;
      17'd68239: data = 8'h04;
      17'd68240: data = 8'h02;
      17'd68241: data = 8'h01;
      17'd68242: data = 8'h02;
      17'd68243: data = 8'h02;
      17'd68244: data = 8'h00;
      17'd68245: data = 8'h00;
      17'd68246: data = 8'h01;
      17'd68247: data = 8'hfd;
      17'd68248: data = 8'hfc;
      17'd68249: data = 8'hfe;
      17'd68250: data = 8'h00;
      17'd68251: data = 8'h00;
      17'd68252: data = 8'h01;
      17'd68253: data = 8'h01;
      17'd68254: data = 8'h00;
      17'd68255: data = 8'h00;
      17'd68256: data = 8'h00;
      17'd68257: data = 8'hfd;
      17'd68258: data = 8'hfd;
      17'd68259: data = 8'hfe;
      17'd68260: data = 8'h01;
      17'd68261: data = 8'h00;
      17'd68262: data = 8'hfd;
      17'd68263: data = 8'hfe;
      17'd68264: data = 8'hfe;
      17'd68265: data = 8'hfd;
      17'd68266: data = 8'hfd;
      17'd68267: data = 8'hfd;
      17'd68268: data = 8'hfe;
      17'd68269: data = 8'h00;
      17'd68270: data = 8'h01;
      17'd68271: data = 8'h02;
      17'd68272: data = 8'h02;
      17'd68273: data = 8'h04;
      17'd68274: data = 8'h02;
      17'd68275: data = 8'h01;
      17'd68276: data = 8'h00;
      17'd68277: data = 8'h00;
      17'd68278: data = 8'h00;
      17'd68279: data = 8'hfd;
      17'd68280: data = 8'h02;
      17'd68281: data = 8'h04;
      17'd68282: data = 8'h02;
      17'd68283: data = 8'h04;
      17'd68284: data = 8'h05;
      17'd68285: data = 8'h04;
      17'd68286: data = 8'h04;
      17'd68287: data = 8'h04;
      17'd68288: data = 8'h04;
      17'd68289: data = 8'h01;
      17'd68290: data = 8'h00;
      17'd68291: data = 8'h01;
      17'd68292: data = 8'h01;
      17'd68293: data = 8'h00;
      17'd68294: data = 8'h00;
      17'd68295: data = 8'h04;
      17'd68296: data = 8'h02;
      17'd68297: data = 8'h02;
      17'd68298: data = 8'h04;
      17'd68299: data = 8'h04;
      17'd68300: data = 8'h04;
      17'd68301: data = 8'h04;
      17'd68302: data = 8'h02;
      17'd68303: data = 8'h00;
      17'd68304: data = 8'h01;
      17'd68305: data = 8'h02;
      17'd68306: data = 8'h01;
      17'd68307: data = 8'h00;
      17'd68308: data = 8'h01;
      17'd68309: data = 8'h01;
      17'd68310: data = 8'h02;
      17'd68311: data = 8'h02;
      17'd68312: data = 8'h01;
      17'd68313: data = 8'h02;
      17'd68314: data = 8'h04;
      17'd68315: data = 8'h01;
      17'd68316: data = 8'h01;
      17'd68317: data = 8'h00;
      17'd68318: data = 8'h01;
      17'd68319: data = 8'h02;
      17'd68320: data = 8'h01;
      17'd68321: data = 8'h01;
      17'd68322: data = 8'h00;
      17'd68323: data = 8'h00;
      17'd68324: data = 8'h00;
      17'd68325: data = 8'h01;
      17'd68326: data = 8'h01;
      17'd68327: data = 8'h02;
      17'd68328: data = 8'h01;
      17'd68329: data = 8'h01;
      17'd68330: data = 8'h00;
      17'd68331: data = 8'hfe;
      17'd68332: data = 8'h00;
      17'd68333: data = 8'hfe;
      17'd68334: data = 8'h00;
      17'd68335: data = 8'h02;
      17'd68336: data = 8'h01;
      17'd68337: data = 8'h01;
      17'd68338: data = 8'h01;
      17'd68339: data = 8'h00;
      17'd68340: data = 8'h00;
      17'd68341: data = 8'h00;
      17'd68342: data = 8'h01;
      17'd68343: data = 8'h00;
      17'd68344: data = 8'h00;
      17'd68345: data = 8'h01;
      17'd68346: data = 8'h01;
      17'd68347: data = 8'h01;
      17'd68348: data = 8'h01;
      17'd68349: data = 8'h01;
      17'd68350: data = 8'h01;
      17'd68351: data = 8'h00;
      17'd68352: data = 8'h00;
      17'd68353: data = 8'h00;
      17'd68354: data = 8'hfe;
      17'd68355: data = 8'hfe;
      17'd68356: data = 8'hfe;
      17'd68357: data = 8'hfe;
      17'd68358: data = 8'h01;
      17'd68359: data = 8'h00;
      17'd68360: data = 8'h00;
      17'd68361: data = 8'h00;
      17'd68362: data = 8'hfe;
      17'd68363: data = 8'hfd;
      17'd68364: data = 8'hfe;
      17'd68365: data = 8'h01;
      17'd68366: data = 8'hfe;
      17'd68367: data = 8'hfd;
      17'd68368: data = 8'hfe;
      17'd68369: data = 8'hfc;
      17'd68370: data = 8'hfc;
      17'd68371: data = 8'hfa;
      17'd68372: data = 8'hfa;
      17'd68373: data = 8'hfa;
      17'd68374: data = 8'hfa;
      17'd68375: data = 8'hf9;
      17'd68376: data = 8'hfa;
      17'd68377: data = 8'hfc;
      17'd68378: data = 8'hfa;
      17'd68379: data = 8'hfc;
      17'd68380: data = 8'hfa;
      17'd68381: data = 8'hf9;
      17'd68382: data = 8'hf9;
      17'd68383: data = 8'hf6;
      17'd68384: data = 8'hf6;
      17'd68385: data = 8'hf5;
      17'd68386: data = 8'hf9;
      17'd68387: data = 8'hfa;
      17'd68388: data = 8'hf9;
      17'd68389: data = 8'hfa;
      17'd68390: data = 8'hf9;
      17'd68391: data = 8'hf9;
      17'd68392: data = 8'hf9;
      17'd68393: data = 8'hf9;
      17'd68394: data = 8'hf6;
      17'd68395: data = 8'hf9;
      17'd68396: data = 8'hf9;
      17'd68397: data = 8'hf6;
      17'd68398: data = 8'hfa;
      17'd68399: data = 8'hfa;
      17'd68400: data = 8'hfa;
      17'd68401: data = 8'hfa;
      17'd68402: data = 8'hf9;
      17'd68403: data = 8'hf6;
      17'd68404: data = 8'hf6;
      17'd68405: data = 8'hf9;
      17'd68406: data = 8'hf9;
      17'd68407: data = 8'hf9;
      17'd68408: data = 8'hfa;
      17'd68409: data = 8'hfa;
      17'd68410: data = 8'hfc;
      17'd68411: data = 8'hfd;
      17'd68412: data = 8'hfc;
      17'd68413: data = 8'hfc;
      17'd68414: data = 8'hf9;
      17'd68415: data = 8'hfa;
      17'd68416: data = 8'hfc;
      17'd68417: data = 8'hfd;
      17'd68418: data = 8'hfc;
      17'd68419: data = 8'hfc;
      17'd68420: data = 8'hfc;
      17'd68421: data = 8'hfc;
      17'd68422: data = 8'hfd;
      17'd68423: data = 8'hfc;
      17'd68424: data = 8'hfc;
      17'd68425: data = 8'hfc;
      17'd68426: data = 8'hfa;
      17'd68427: data = 8'hfc;
      17'd68428: data = 8'hfc;
      17'd68429: data = 8'hfa;
      17'd68430: data = 8'hfa;
      17'd68431: data = 8'hfc;
      17'd68432: data = 8'hfc;
      17'd68433: data = 8'hfa;
      17'd68434: data = 8'hf9;
      17'd68435: data = 8'hfc;
      17'd68436: data = 8'hfc;
      17'd68437: data = 8'hfc;
      17'd68438: data = 8'hfc;
      17'd68439: data = 8'hfc;
      17'd68440: data = 8'hfd;
      17'd68441: data = 8'hfd;
      17'd68442: data = 8'hfe;
      17'd68443: data = 8'hfd;
      17'd68444: data = 8'hfc;
      17'd68445: data = 8'hfc;
      17'd68446: data = 8'hfc;
      17'd68447: data = 8'hfc;
      17'd68448: data = 8'hfc;
      17'd68449: data = 8'hfd;
      17'd68450: data = 8'hfd;
      17'd68451: data = 8'hfe;
      17'd68452: data = 8'hfd;
      17'd68453: data = 8'h00;
      17'd68454: data = 8'h00;
      17'd68455: data = 8'h06;
      17'd68456: data = 8'h09;
      17'd68457: data = 8'hf6;
      17'd68458: data = 8'hf6;
      17'd68459: data = 8'hec;
      17'd68460: data = 8'heb;
      17'd68461: data = 8'hf4;
      17'd68462: data = 8'h00;
      17'd68463: data = 8'h0c;
      17'd68464: data = 8'h1b;
      17'd68465: data = 8'h23;
      17'd68466: data = 8'h1f;
      17'd68467: data = 8'h0e;
      17'd68468: data = 8'hf4;
      17'd68469: data = 8'he4;
      17'd68470: data = 8'hd6;
      17'd68471: data = 8'he0;
      17'd68472: data = 8'hf6;
      17'd68473: data = 8'h0d;
      17'd68474: data = 8'h1f;
      17'd68475: data = 8'h29;
      17'd68476: data = 8'h24;
      17'd68477: data = 8'h15;
      17'd68478: data = 8'h09;
      17'd68479: data = 8'hfd;
      17'd68480: data = 8'hf4;
      17'd68481: data = 8'hfc;
      17'd68482: data = 8'h01;
      17'd68483: data = 8'h02;
      17'd68484: data = 8'h04;
      17'd68485: data = 8'hfd;
      17'd68486: data = 8'hfa;
      17'd68487: data = 8'hfa;
      17'd68488: data = 8'hf2;
      17'd68489: data = 8'hf9;
      17'd68490: data = 8'h05;
      17'd68491: data = 8'h0a;
      17'd68492: data = 8'h0e;
      17'd68493: data = 8'h0d;
      17'd68494: data = 8'h0a;
      17'd68495: data = 8'h04;
      17'd68496: data = 8'hf4;
      17'd68497: data = 8'he9;
      17'd68498: data = 8'hec;
      17'd68499: data = 8'hf6;
      17'd68500: data = 8'hfe;
      17'd68501: data = 8'h04;
      17'd68502: data = 8'h06;
      17'd68503: data = 8'h06;
      17'd68504: data = 8'h02;
      17'd68505: data = 8'hfc;
      17'd68506: data = 8'h02;
      17'd68507: data = 8'h05;
      17'd68508: data = 8'hfd;
      17'd68509: data = 8'h02;
      17'd68510: data = 8'h0a;
      17'd68511: data = 8'h0a;
      17'd68512: data = 8'h02;
      17'd68513: data = 8'hfe;
      17'd68514: data = 8'h00;
      17'd68515: data = 8'h00;
      17'd68516: data = 8'h01;
      17'd68517: data = 8'h06;
      17'd68518: data = 8'h0a;
      17'd68519: data = 8'h0e;
      17'd68520: data = 8'h0d;
      17'd68521: data = 8'h06;
      17'd68522: data = 8'h06;
      17'd68523: data = 8'h0c;
      17'd68524: data = 8'h0e;
      17'd68525: data = 8'h0e;
      17'd68526: data = 8'h12;
      17'd68527: data = 8'h15;
      17'd68528: data = 8'h11;
      17'd68529: data = 8'h05;
      17'd68530: data = 8'h01;
      17'd68531: data = 8'hfe;
      17'd68532: data = 8'h00;
      17'd68533: data = 8'h09;
      17'd68534: data = 8'h0a;
      17'd68535: data = 8'h09;
      17'd68536: data = 8'h0e;
      17'd68537: data = 8'h12;
      17'd68538: data = 8'h12;
      17'd68539: data = 8'h0e;
      17'd68540: data = 8'h0a;
      17'd68541: data = 8'h01;
      17'd68542: data = 8'hfe;
      17'd68543: data = 8'h04;
      17'd68544: data = 8'h04;
      17'd68545: data = 8'h06;
      17'd68546: data = 8'h0a;
      17'd68547: data = 8'h05;
      17'd68548: data = 8'hfe;
      17'd68549: data = 8'hf9;
      17'd68550: data = 8'hf2;
      17'd68551: data = 8'hf4;
      17'd68552: data = 8'hfe;
      17'd68553: data = 8'h06;
      17'd68554: data = 8'h0a;
      17'd68555: data = 8'h09;
      17'd68556: data = 8'h0a;
      17'd68557: data = 8'hfd;
      17'd68558: data = 8'hf5;
      17'd68559: data = 8'hf4;
      17'd68560: data = 8'hf4;
      17'd68561: data = 8'h00;
      17'd68562: data = 8'h05;
      17'd68563: data = 8'hfe;
      17'd68564: data = 8'hf4;
      17'd68565: data = 8'hf2;
      17'd68566: data = 8'hf6;
      17'd68567: data = 8'hfd;
      17'd68568: data = 8'h01;
      17'd68569: data = 8'h04;
      17'd68570: data = 8'hfe;
      17'd68571: data = 8'hf9;
      17'd68572: data = 8'hfa;
      17'd68573: data = 8'hfd;
      17'd68574: data = 8'hfd;
      17'd68575: data = 8'h02;
      17'd68576: data = 8'h02;
      17'd68577: data = 8'hfc;
      17'd68578: data = 8'hf5;
      17'd68579: data = 8'heb;
      17'd68580: data = 8'hef;
      17'd68581: data = 8'hfa;
      17'd68582: data = 8'hfe;
      17'd68583: data = 8'hfd;
      17'd68584: data = 8'h00;
      17'd68585: data = 8'h04;
      17'd68586: data = 8'h00;
      17'd68587: data = 8'hfa;
      17'd68588: data = 8'hfc;
      17'd68589: data = 8'hfd;
      17'd68590: data = 8'hfe;
      17'd68591: data = 8'hfe;
      17'd68592: data = 8'hf9;
      17'd68593: data = 8'hf5;
      17'd68594: data = 8'hf4;
      17'd68595: data = 8'hf5;
      17'd68596: data = 8'hfd;
      17'd68597: data = 8'hfe;
      17'd68598: data = 8'hfc;
      17'd68599: data = 8'hf6;
      17'd68600: data = 8'hf6;
      17'd68601: data = 8'hfc;
      17'd68602: data = 8'h01;
      17'd68603: data = 8'h01;
      17'd68604: data = 8'h00;
      17'd68605: data = 8'h00;
      17'd68606: data = 8'hfe;
      17'd68607: data = 8'hfa;
      17'd68608: data = 8'hf5;
      17'd68609: data = 8'hfa;
      17'd68610: data = 8'hfc;
      17'd68611: data = 8'hfc;
      17'd68612: data = 8'h01;
      17'd68613: data = 8'h01;
      17'd68614: data = 8'hfe;
      17'd68615: data = 8'hfd;
      17'd68616: data = 8'hf6;
      17'd68617: data = 8'hfd;
      17'd68618: data = 8'h06;
      17'd68619: data = 8'h02;
      17'd68620: data = 8'hfe;
      17'd68621: data = 8'h00;
      17'd68622: data = 8'h01;
      17'd68623: data = 8'hfe;
      17'd68624: data = 8'hf6;
      17'd68625: data = 8'hfa;
      17'd68626: data = 8'hf9;
      17'd68627: data = 8'hfa;
      17'd68628: data = 8'hfd;
      17'd68629: data = 8'h02;
      17'd68630: data = 8'h0a;
      17'd68631: data = 8'h0c;
      17'd68632: data = 8'h04;
      17'd68633: data = 8'h05;
      17'd68634: data = 8'h00;
      17'd68635: data = 8'hfc;
      17'd68636: data = 8'h05;
      17'd68637: data = 8'h0a;
      17'd68638: data = 8'h0c;
      17'd68639: data = 8'h04;
      17'd68640: data = 8'hfe;
      17'd68641: data = 8'hfe;
      17'd68642: data = 8'hf9;
      17'd68643: data = 8'hf6;
      17'd68644: data = 8'h04;
      17'd68645: data = 8'h06;
      17'd68646: data = 8'h04;
      17'd68647: data = 8'h0a;
      17'd68648: data = 8'h05;
      17'd68649: data = 8'hfe;
      17'd68650: data = 8'hfd;
      17'd68651: data = 8'hf9;
      17'd68652: data = 8'hf9;
      17'd68653: data = 8'hfd;
      17'd68654: data = 8'h00;
      17'd68655: data = 8'h00;
      17'd68656: data = 8'hfe;
      17'd68657: data = 8'hfe;
      17'd68658: data = 8'hfe;
      17'd68659: data = 8'hfd;
      17'd68660: data = 8'h00;
      17'd68661: data = 8'h01;
      17'd68662: data = 8'h05;
      17'd68663: data = 8'h04;
      17'd68664: data = 8'hfe;
      17'd68665: data = 8'hfa;
      17'd68666: data = 8'hfe;
      17'd68667: data = 8'h02;
      17'd68668: data = 8'h02;
      17'd68669: data = 8'h05;
      17'd68670: data = 8'h01;
      17'd68671: data = 8'hfd;
      17'd68672: data = 8'hfd;
      17'd68673: data = 8'h01;
      17'd68674: data = 8'h04;
      17'd68675: data = 8'h06;
      17'd68676: data = 8'h09;
      17'd68677: data = 8'h0d;
      17'd68678: data = 8'h0c;
      17'd68679: data = 8'h06;
      17'd68680: data = 8'h04;
      17'd68681: data = 8'h04;
      17'd68682: data = 8'h09;
      17'd68683: data = 8'h0d;
      17'd68684: data = 8'h06;
      17'd68685: data = 8'h04;
      17'd68686: data = 8'h02;
      17'd68687: data = 8'h01;
      17'd68688: data = 8'h00;
      17'd68689: data = 8'h00;
      17'd68690: data = 8'h04;
      17'd68691: data = 8'h09;
      17'd68692: data = 8'h05;
      17'd68693: data = 8'h09;
      17'd68694: data = 8'h0a;
      17'd68695: data = 8'h05;
      17'd68696: data = 8'h01;
      17'd68697: data = 8'h02;
      17'd68698: data = 8'h04;
      17'd68699: data = 8'h00;
      17'd68700: data = 8'hfd;
      17'd68701: data = 8'hfd;
      17'd68702: data = 8'hfa;
      17'd68703: data = 8'hf9;
      17'd68704: data = 8'hf6;
      17'd68705: data = 8'hf6;
      17'd68706: data = 8'hfc;
      17'd68707: data = 8'h00;
      17'd68708: data = 8'hfc;
      17'd68709: data = 8'hf9;
      17'd68710: data = 8'hfd;
      17'd68711: data = 8'hfc;
      17'd68712: data = 8'hfd;
      17'd68713: data = 8'hfc;
      17'd68714: data = 8'hfc;
      17'd68715: data = 8'hf5;
      17'd68716: data = 8'hf4;
      17'd68717: data = 8'hf2;
      17'd68718: data = 8'hef;
      17'd68719: data = 8'hf5;
      17'd68720: data = 8'hf4;
      17'd68721: data = 8'hf9;
      17'd68722: data = 8'hfd;
      17'd68723: data = 8'hfd;
      17'd68724: data = 8'hfe;
      17'd68725: data = 8'hfc;
      17'd68726: data = 8'hf5;
      17'd68727: data = 8'hfd;
      17'd68728: data = 8'hfe;
      17'd68729: data = 8'h00;
      17'd68730: data = 8'h02;
      17'd68731: data = 8'hf6;
      17'd68732: data = 8'hf9;
      17'd68733: data = 8'hf6;
      17'd68734: data = 8'hf4;
      17'd68735: data = 8'h00;
      17'd68736: data = 8'hfd;
      17'd68737: data = 8'hfe;
      17'd68738: data = 8'h06;
      17'd68739: data = 8'h02;
      17'd68740: data = 8'h01;
      17'd68741: data = 8'h06;
      17'd68742: data = 8'hfc;
      17'd68743: data = 8'h02;
      17'd68744: data = 8'h02;
      17'd68745: data = 8'hf9;
      17'd68746: data = 8'hfd;
      17'd68747: data = 8'hf6;
      17'd68748: data = 8'hef;
      17'd68749: data = 8'hf5;
      17'd68750: data = 8'hec;
      17'd68751: data = 8'hf2;
      17'd68752: data = 8'h00;
      17'd68753: data = 8'h00;
      17'd68754: data = 8'h09;
      17'd68755: data = 8'h09;
      17'd68756: data = 8'hfc;
      17'd68757: data = 8'h02;
      17'd68758: data = 8'hfd;
      17'd68759: data = 8'h02;
      17'd68760: data = 8'h0d;
      17'd68761: data = 8'h04;
      17'd68762: data = 8'h06;
      17'd68763: data = 8'hfc;
      17'd68764: data = 8'hf2;
      17'd68765: data = 8'hf9;
      17'd68766: data = 8'hfc;
      17'd68767: data = 8'h04;
      17'd68768: data = 8'h13;
      17'd68769: data = 8'h0d;
      17'd68770: data = 8'h06;
      17'd68771: data = 8'h04;
      17'd68772: data = 8'hfd;
      17'd68773: data = 8'h09;
      17'd68774: data = 8'h0e;
      17'd68775: data = 8'h11;
      17'd68776: data = 8'h0d;
      17'd68777: data = 8'h00;
      17'd68778: data = 8'hf1;
      17'd68779: data = 8'hec;
      17'd68780: data = 8'hed;
      17'd68781: data = 8'hf5;
      17'd68782: data = 8'hfd;
      17'd68783: data = 8'hfc;
      17'd68784: data = 8'hf6;
      17'd68785: data = 8'hed;
      17'd68786: data = 8'heb;
      17'd68787: data = 8'heb;
      17'd68788: data = 8'hf4;
      17'd68789: data = 8'hf9;
      17'd68790: data = 8'hf9;
      17'd68791: data = 8'hf2;
      17'd68792: data = 8'he3;
      17'd68793: data = 8'hdb;
      17'd68794: data = 8'hd8;
      17'd68795: data = 8'hdc;
      17'd68796: data = 8'he7;
      17'd68797: data = 8'hec;
      17'd68798: data = 8'heb;
      17'd68799: data = 8'he5;
      17'd68800: data = 8'he0;
      17'd68801: data = 8'he4;
      17'd68802: data = 8'hef;
      17'd68803: data = 8'hf5;
      17'd68804: data = 8'h04;
      17'd68805: data = 8'h04;
      17'd68806: data = 8'hfd;
      17'd68807: data = 8'hf9;
      17'd68808: data = 8'hf4;
      17'd68809: data = 8'hfc;
      17'd68810: data = 8'h04;
      17'd68811: data = 8'h09;
      17'd68812: data = 8'h0d;
      17'd68813: data = 8'h0c;
      17'd68814: data = 8'h09;
      17'd68815: data = 8'h09;
      17'd68816: data = 8'h0d;
      17'd68817: data = 8'h1f;
      17'd68818: data = 8'h27;
      17'd68819: data = 8'h29;
      17'd68820: data = 8'h29;
      17'd68821: data = 8'h1e;
      17'd68822: data = 8'h1a;
      17'd68823: data = 8'h1b;
      17'd68824: data = 8'h1c;
      17'd68825: data = 8'h23;
      17'd68826: data = 8'h26;
      17'd68827: data = 8'h1c;
      17'd68828: data = 8'h19;
      17'd68829: data = 8'h13;
      17'd68830: data = 8'h13;
      17'd68831: data = 8'h19;
      17'd68832: data = 8'h1b;
      17'd68833: data = 8'h1e;
      17'd68834: data = 8'h1a;
      17'd68835: data = 8'h11;
      17'd68836: data = 8'h0c;
      17'd68837: data = 8'h05;
      17'd68838: data = 8'h06;
      17'd68839: data = 8'h06;
      17'd68840: data = 8'h02;
      17'd68841: data = 8'hfe;
      17'd68842: data = 8'hf4;
      17'd68843: data = 8'hec;
      17'd68844: data = 8'heb;
      17'd68845: data = 8'hec;
      17'd68846: data = 8'hf2;
      17'd68847: data = 8'hf4;
      17'd68848: data = 8'hf1;
      17'd68849: data = 8'hed;
      17'd68850: data = 8'hec;
      17'd68851: data = 8'he9;
      17'd68852: data = 8'he9;
      17'd68853: data = 8'hef;
      17'd68854: data = 8'hf1;
      17'd68855: data = 8'hef;
      17'd68856: data = 8'hef;
      17'd68857: data = 8'hec;
      17'd68858: data = 8'he9;
      17'd68859: data = 8'hec;
      17'd68860: data = 8'hed;
      17'd68861: data = 8'hf4;
      17'd68862: data = 8'hfa;
      17'd68863: data = 8'hfd;
      17'd68864: data = 8'h01;
      17'd68865: data = 8'h02;
      17'd68866: data = 8'h01;
      17'd68867: data = 8'h01;
      17'd68868: data = 8'h01;
      17'd68869: data = 8'h04;
      17'd68870: data = 8'h0c;
      17'd68871: data = 8'h12;
      17'd68872: data = 8'h16;
      17'd68873: data = 8'h15;
      17'd68874: data = 8'h0c;
      17'd68875: data = 8'h09;
      17'd68876: data = 8'h09;
      17'd68877: data = 8'h0c;
      17'd68878: data = 8'h12;
      17'd68879: data = 8'h19;
      17'd68880: data = 8'h15;
      17'd68881: data = 8'h0e;
      17'd68882: data = 8'h06;
      17'd68883: data = 8'h04;
      17'd68884: data = 8'h06;
      17'd68885: data = 8'h0a;
      17'd68886: data = 8'h0d;
      17'd68887: data = 8'h0a;
      17'd68888: data = 8'h01;
      17'd68889: data = 8'hfc;
      17'd68890: data = 8'hf9;
      17'd68891: data = 8'hf9;
      17'd68892: data = 8'hfc;
      17'd68893: data = 8'hf9;
      17'd68894: data = 8'hf2;
      17'd68895: data = 8'he9;
      17'd68896: data = 8'he4;
      17'd68897: data = 8'he5;
      17'd68898: data = 8'hec;
      17'd68899: data = 8'hef;
      17'd68900: data = 8'hef;
      17'd68901: data = 8'hef;
      17'd68902: data = 8'he5;
      17'd68903: data = 8'he0;
      17'd68904: data = 8'hde;
      17'd68905: data = 8'he0;
      17'd68906: data = 8'he5;
      17'd68907: data = 8'he9;
      17'd68908: data = 8'heb;
      17'd68909: data = 8'he7;
      17'd68910: data = 8'he5;
      17'd68911: data = 8'he5;
      17'd68912: data = 8'he7;
      17'd68913: data = 8'heb;
      17'd68914: data = 8'hf1;
      17'd68915: data = 8'hf9;
      17'd68916: data = 8'hfc;
      17'd68917: data = 8'hfa;
      17'd68918: data = 8'h00;
      17'd68919: data = 8'h00;
      17'd68920: data = 8'h01;
      17'd68921: data = 8'h06;
      17'd68922: data = 8'h04;
      17'd68923: data = 8'h06;
      17'd68924: data = 8'h09;
      17'd68925: data = 8'h04;
      17'd68926: data = 8'h0e;
      17'd68927: data = 8'h0d;
      17'd68928: data = 8'h11;
      17'd68929: data = 8'h16;
      17'd68930: data = 8'h11;
      17'd68931: data = 8'h12;
      17'd68932: data = 8'h0e;
      17'd68933: data = 8'h0c;
      17'd68934: data = 8'h12;
      17'd68935: data = 8'h0e;
      17'd68936: data = 8'h12;
      17'd68937: data = 8'h15;
      17'd68938: data = 8'h0d;
      17'd68939: data = 8'h0c;
      17'd68940: data = 8'h06;
      17'd68941: data = 8'h01;
      17'd68942: data = 8'h00;
      17'd68943: data = 8'h00;
      17'd68944: data = 8'h00;
      17'd68945: data = 8'hfd;
      17'd68946: data = 8'h00;
      17'd68947: data = 8'hfc;
      17'd68948: data = 8'hf9;
      17'd68949: data = 8'hfd;
      17'd68950: data = 8'hf5;
      17'd68951: data = 8'hf9;
      17'd68952: data = 8'hfe;
      17'd68953: data = 8'hf6;
      17'd68954: data = 8'hfc;
      17'd68955: data = 8'hf5;
      17'd68956: data = 8'hf5;
      17'd68957: data = 8'hf6;
      17'd68958: data = 8'hf9;
      17'd68959: data = 8'hf6;
      17'd68960: data = 8'hf9;
      17'd68961: data = 8'hf9;
      17'd68962: data = 8'h01;
      17'd68963: data = 8'h01;
      17'd68964: data = 8'h06;
      17'd68965: data = 8'h05;
      17'd68966: data = 8'h05;
      17'd68967: data = 8'h06;
      17'd68968: data = 8'h04;
      17'd68969: data = 8'h06;
      17'd68970: data = 8'h13;
      17'd68971: data = 8'h11;
      17'd68972: data = 8'h0a;
      17'd68973: data = 8'h15;
      17'd68974: data = 8'h06;
      17'd68975: data = 8'h09;
      17'd68976: data = 8'h0d;
      17'd68977: data = 8'h06;
      17'd68978: data = 8'h12;
      17'd68979: data = 8'h15;
      17'd68980: data = 8'h0a;
      17'd68981: data = 8'h1c;
      17'd68982: data = 8'h1c;
      17'd68983: data = 8'h15;
      17'd68984: data = 8'h1a;
      17'd68985: data = 8'h0a;
      17'd68986: data = 8'h01;
      17'd68987: data = 8'h04;
      17'd68988: data = 8'h01;
      17'd68989: data = 8'h02;
      17'd68990: data = 8'h04;
      17'd68991: data = 8'h01;
      17'd68992: data = 8'hfc;
      17'd68993: data = 8'hfa;
      17'd68994: data = 8'hf2;
      17'd68995: data = 8'hf6;
      17'd68996: data = 8'h04;
      17'd68997: data = 8'h0c;
      17'd68998: data = 8'h12;
      17'd68999: data = 8'h19;
      17'd69000: data = 8'h13;
      17'd69001: data = 8'h11;
      17'd69002: data = 8'h0a;
      17'd69003: data = 8'h0d;
      17'd69004: data = 8'h0e;
      17'd69005: data = 8'h06;
      17'd69006: data = 8'h0d;
      17'd69007: data = 8'h09;
      17'd69008: data = 8'h02;
      17'd69009: data = 8'h0a;
      17'd69010: data = 8'h05;
      17'd69011: data = 8'h0d;
      17'd69012: data = 8'h0e;
      17'd69013: data = 8'h06;
      17'd69014: data = 8'h0a;
      17'd69015: data = 8'h05;
      17'd69016: data = 8'hfe;
      17'd69017: data = 8'h06;
      17'd69018: data = 8'h06;
      17'd69019: data = 8'h04;
      17'd69020: data = 8'h01;
      17'd69021: data = 8'hf1;
      17'd69022: data = 8'he9;
      17'd69023: data = 8'hdb;
      17'd69024: data = 8'hdb;
      17'd69025: data = 8'he0;
      17'd69026: data = 8'he0;
      17'd69027: data = 8'he5;
      17'd69028: data = 8'he0;
      17'd69029: data = 8'hda;
      17'd69030: data = 8'hd5;
      17'd69031: data = 8'hce;
      17'd69032: data = 8'hd5;
      17'd69033: data = 8'hd6;
      17'd69034: data = 8'hd6;
      17'd69035: data = 8'hde;
      17'd69036: data = 8'hd6;
      17'd69037: data = 8'hd2;
      17'd69038: data = 8'hcd;
      17'd69039: data = 8'hcd;
      17'd69040: data = 8'hd1;
      17'd69041: data = 8'hd1;
      17'd69042: data = 8'hd8;
      17'd69043: data = 8'hdc;
      17'd69044: data = 8'hde;
      17'd69045: data = 8'he5;
      17'd69046: data = 8'hef;
      17'd69047: data = 8'hfa;
      17'd69048: data = 8'h06;
      17'd69049: data = 8'h0c;
      17'd69050: data = 8'h11;
      17'd69051: data = 8'h13;
      17'd69052: data = 8'h11;
      17'd69053: data = 8'h15;
      17'd69054: data = 8'h1e;
      17'd69055: data = 8'h22;
      17'd69056: data = 8'h24;
      17'd69057: data = 8'h24;
      17'd69058: data = 8'h23;
      17'd69059: data = 8'h22;
      17'd69060: data = 8'h27;
      17'd69061: data = 8'h2d;
      17'd69062: data = 8'h31;
      17'd69063: data = 8'h35;
      17'd69064: data = 8'h36;
      17'd69065: data = 8'h33;
      17'd69066: data = 8'h31;
      17'd69067: data = 8'h2c;
      17'd69068: data = 8'h24;
      17'd69069: data = 8'h23;
      17'd69070: data = 8'h19;
      17'd69071: data = 8'h0e;
      17'd69072: data = 8'h0c;
      17'd69073: data = 8'h00;
      17'd69074: data = 8'hfa;
      17'd69075: data = 8'hf6;
      17'd69076: data = 8'hf4;
      17'd69077: data = 8'hef;
      17'd69078: data = 8'hef;
      17'd69079: data = 8'heb;
      17'd69080: data = 8'he7;
      17'd69081: data = 8'he3;
      17'd69082: data = 8'he2;
      17'd69083: data = 8'hde;
      17'd69084: data = 8'hdc;
      17'd69085: data = 8'hdb;
      17'd69086: data = 8'hd5;
      17'd69087: data = 8'hd2;
      17'd69088: data = 8'hcb;
      17'd69089: data = 8'hcb;
      17'd69090: data = 8'hcb;
      17'd69091: data = 8'hce;
      17'd69092: data = 8'hd6;
      17'd69093: data = 8'he0;
      17'd69094: data = 8'he5;
      17'd69095: data = 8'heb;
      17'd69096: data = 8'hf1;
      17'd69097: data = 8'hf9;
      17'd69098: data = 8'h00;
      17'd69099: data = 8'h05;
      17'd69100: data = 8'h0c;
      17'd69101: data = 8'h0d;
      17'd69102: data = 8'h0e;
      17'd69103: data = 8'h0e;
      17'd69104: data = 8'h12;
      17'd69105: data = 8'h15;
      17'd69106: data = 8'h16;
      17'd69107: data = 8'h1a;
      17'd69108: data = 8'h1e;
      17'd69109: data = 8'h1f;
      17'd69110: data = 8'h1f;
      17'd69111: data = 8'h22;
      17'd69112: data = 8'h26;
      17'd69113: data = 8'h29;
      17'd69114: data = 8'h29;
      17'd69115: data = 8'h29;
      17'd69116: data = 8'h24;
      17'd69117: data = 8'h1b;
      17'd69118: data = 8'h13;
      17'd69119: data = 8'h0a;
      17'd69120: data = 8'h05;
      17'd69121: data = 8'h01;
      17'd69122: data = 8'hfd;
      17'd69123: data = 8'hf6;
      17'd69124: data = 8'hec;
      17'd69125: data = 8'he4;
      17'd69126: data = 8'he2;
      17'd69127: data = 8'hdc;
      17'd69128: data = 8'he0;
      17'd69129: data = 8'he4;
      17'd69130: data = 8'he4;
      17'd69131: data = 8'he5;
      17'd69132: data = 8'hda;
      17'd69133: data = 8'hd2;
      17'd69134: data = 8'hd1;
      17'd69135: data = 8'hc6;
      17'd69136: data = 8'hcb;
      17'd69137: data = 8'hcb;
      17'd69138: data = 8'hc9;
      17'd69139: data = 8'hcb;
      17'd69140: data = 8'hcb;
      17'd69141: data = 8'hd3;
      17'd69142: data = 8'hde;
      17'd69143: data = 8'he5;
      17'd69144: data = 8'hf1;
      17'd69145: data = 8'hf1;
      17'd69146: data = 8'hf6;
      17'd69147: data = 8'hfd;
      17'd69148: data = 8'h02;
      17'd69149: data = 8'h12;
      17'd69150: data = 8'h15;
      17'd69151: data = 8'h15;
      17'd69152: data = 8'h16;
      17'd69153: data = 8'h0e;
      17'd69154: data = 8'h0e;
      17'd69155: data = 8'h13;
      17'd69156: data = 8'h19;
      17'd69157: data = 8'h26;
      17'd69158: data = 8'h2b;
      17'd69159: data = 8'h31;
      17'd69160: data = 8'h34;
      17'd69161: data = 8'h33;
      17'd69162: data = 8'h34;
      17'd69163: data = 8'h2d;
      17'd69164: data = 8'h29;
      17'd69165: data = 8'h29;
      17'd69166: data = 8'h1c;
      17'd69167: data = 8'h1a;
      17'd69168: data = 8'h15;
      17'd69169: data = 8'h0c;
      17'd69170: data = 8'h0c;
      17'd69171: data = 8'h01;
      17'd69172: data = 8'hfc;
      17'd69173: data = 8'hfa;
      17'd69174: data = 8'hf1;
      17'd69175: data = 8'hf1;
      17'd69176: data = 8'hf2;
      17'd69177: data = 8'hf1;
      17'd69178: data = 8'hf6;
      17'd69179: data = 8'hf2;
      17'd69180: data = 8'he9;
      17'd69181: data = 8'he5;
      17'd69182: data = 8'hdc;
      17'd69183: data = 8'hdc;
      17'd69184: data = 8'he0;
      17'd69185: data = 8'hdc;
      17'd69186: data = 8'hde;
      17'd69187: data = 8'he3;
      17'd69188: data = 8'he2;
      17'd69189: data = 8'he7;
      17'd69190: data = 8'hef;
      17'd69191: data = 8'hf1;
      17'd69192: data = 8'hfd;
      17'd69193: data = 8'h01;
      17'd69194: data = 8'h02;
      17'd69195: data = 8'h0d;
      17'd69196: data = 8'h0d;
      17'd69197: data = 8'h0e;
      17'd69198: data = 8'h13;
      17'd69199: data = 8'h11;
      17'd69200: data = 8'h0e;
      17'd69201: data = 8'h11;
      17'd69202: data = 8'h0d;
      17'd69203: data = 8'h15;
      17'd69204: data = 8'h1b;
      17'd69205: data = 8'h1f;
      17'd69206: data = 8'h23;
      17'd69207: data = 8'h19;
      17'd69208: data = 8'h1b;
      17'd69209: data = 8'h1e;
      17'd69210: data = 8'h1b;
      17'd69211: data = 8'h23;
      17'd69212: data = 8'h23;
      17'd69213: data = 8'h24;
      17'd69214: data = 8'h26;
      17'd69215: data = 8'h1b;
      17'd69216: data = 8'h1b;
      17'd69217: data = 8'h0d;
      17'd69218: data = 8'h04;
      17'd69219: data = 8'h06;
      17'd69220: data = 8'hf9;
      17'd69221: data = 8'h00;
      17'd69222: data = 8'hfd;
      17'd69223: data = 8'hfc;
      17'd69224: data = 8'h0d;
      17'd69225: data = 8'hfa;
      17'd69226: data = 8'h04;
      17'd69227: data = 8'h11;
      17'd69228: data = 8'hf6;
      17'd69229: data = 8'h0d;
      17'd69230: data = 8'hfc;
      17'd69231: data = 8'hf4;
      17'd69232: data = 8'h05;
      17'd69233: data = 8'hf1;
      17'd69234: data = 8'hef;
      17'd69235: data = 8'hfa;
      17'd69236: data = 8'he0;
      17'd69237: data = 8'hf2;
      17'd69238: data = 8'hf4;
      17'd69239: data = 8'hf5;
      17'd69240: data = 8'h04;
      17'd69241: data = 8'h00;
      17'd69242: data = 8'h02;
      17'd69243: data = 8'h13;
      17'd69244: data = 8'h13;
      17'd69245: data = 8'h11;
      17'd69246: data = 8'h16;
      17'd69247: data = 8'h04;
      17'd69248: data = 8'h04;
      17'd69249: data = 8'hfc;
      17'd69250: data = 8'hf9;
      17'd69251: data = 8'hfa;
      17'd69252: data = 8'h04;
      17'd69253: data = 8'h0e;
      17'd69254: data = 8'h19;
      17'd69255: data = 8'h16;
      17'd69256: data = 8'h1b;
      17'd69257: data = 8'h1b;
      17'd69258: data = 8'h24;
      17'd69259: data = 8'h23;
      17'd69260: data = 8'h29;
      17'd69261: data = 8'h2d;
      17'd69262: data = 8'h27;
      17'd69263: data = 8'h27;
      17'd69264: data = 8'h1c;
      17'd69265: data = 8'h16;
      17'd69266: data = 8'h0c;
      17'd69267: data = 8'h00;
      17'd69268: data = 8'hfe;
      17'd69269: data = 8'hf4;
      17'd69270: data = 8'hf5;
      17'd69271: data = 8'hf9;
      17'd69272: data = 8'hf6;
      17'd69273: data = 8'hfa;
      17'd69274: data = 8'hfd;
      17'd69275: data = 8'hf5;
      17'd69276: data = 8'hf1;
      17'd69277: data = 8'he5;
      17'd69278: data = 8'he3;
      17'd69279: data = 8'hdc;
      17'd69280: data = 8'hd2;
      17'd69281: data = 8'hcd;
      17'd69282: data = 8'hcb;
      17'd69283: data = 8'hc2;
      17'd69284: data = 8'hbb;
      17'd69285: data = 8'hb8;
      17'd69286: data = 8'hb3;
      17'd69287: data = 8'hb5;
      17'd69288: data = 8'hb8;
      17'd69289: data = 8'hc0;
      17'd69290: data = 8'hc6;
      17'd69291: data = 8'hd3;
      17'd69292: data = 8'hdb;
      17'd69293: data = 8'he3;
      17'd69294: data = 8'he2;
      17'd69295: data = 8'hde;
      17'd69296: data = 8'hde;
      17'd69297: data = 8'he0;
      17'd69298: data = 8'he0;
      17'd69299: data = 8'he9;
      17'd69300: data = 8'hed;
      17'd69301: data = 8'hf4;
      17'd69302: data = 8'hf6;
      17'd69303: data = 8'hfe;
      17'd69304: data = 8'h0a;
      17'd69305: data = 8'h0d;
      17'd69306: data = 8'h1a;
      17'd69307: data = 8'h23;
      17'd69308: data = 8'h29;
      17'd69309: data = 8'h33;
      17'd69310: data = 8'h36;
      17'd69311: data = 8'h3d;
      17'd69312: data = 8'h3c;
      17'd69313: data = 8'h39;
      17'd69314: data = 8'h33;
      17'd69315: data = 8'h27;
      17'd69316: data = 8'h1e;
      17'd69317: data = 8'h1c;
      17'd69318: data = 8'h19;
      17'd69319: data = 8'h1b;
      17'd69320: data = 8'h1b;
      17'd69321: data = 8'h1a;
      17'd69322: data = 8'h15;
      17'd69323: data = 8'h0e;
      17'd69324: data = 8'h0a;
      17'd69325: data = 8'h05;
      17'd69326: data = 8'h01;
      17'd69327: data = 8'hfe;
      17'd69328: data = 8'hfc;
      17'd69329: data = 8'hf2;
      17'd69330: data = 8'hec;
      17'd69331: data = 8'he3;
      17'd69332: data = 8'hda;
      17'd69333: data = 8'hd2;
      17'd69334: data = 8'hca;
      17'd69335: data = 8'hc6;
      17'd69336: data = 8'hc9;
      17'd69337: data = 8'hc9;
      17'd69338: data = 8'hce;
      17'd69339: data = 8'hd6;
      17'd69340: data = 8'hde;
      17'd69341: data = 8'he4;
      17'd69342: data = 8'he7;
      17'd69343: data = 8'heb;
      17'd69344: data = 8'heb;
      17'd69345: data = 8'heb;
      17'd69346: data = 8'hed;
      17'd69347: data = 8'hf4;
      17'd69348: data = 8'hf9;
      17'd69349: data = 8'hfe;
      17'd69350: data = 8'hfd;
      17'd69351: data = 8'h01;
      17'd69352: data = 8'h04;
      17'd69353: data = 8'h09;
      17'd69354: data = 8'h11;
      17'd69355: data = 8'h16;
      17'd69356: data = 8'h1e;
      17'd69357: data = 8'h26;
      17'd69358: data = 8'h2b;
      17'd69359: data = 8'h2d;
      17'd69360: data = 8'h2f;
      17'd69361: data = 8'h2c;
      17'd69362: data = 8'h27;
      17'd69363: data = 8'h22;
      17'd69364: data = 8'h1a;
      17'd69365: data = 8'h1a;
      17'd69366: data = 8'h11;
      17'd69367: data = 8'h0a;
      17'd69368: data = 8'h06;
      17'd69369: data = 8'h04;
      17'd69370: data = 8'h00;
      17'd69371: data = 8'hfc;
      17'd69372: data = 8'hf6;
      17'd69373: data = 8'hf5;
      17'd69374: data = 8'hf2;
      17'd69375: data = 8'hf2;
      17'd69376: data = 8'hf4;
      17'd69377: data = 8'hed;
      17'd69378: data = 8'heb;
      17'd69379: data = 8'he4;
      17'd69380: data = 8'hdc;
      17'd69381: data = 8'hda;
      17'd69382: data = 8'hd5;
      17'd69383: data = 8'hd1;
      17'd69384: data = 8'hce;
      17'd69385: data = 8'hd1;
      17'd69386: data = 8'hd8;
      17'd69387: data = 8'hdb;
      17'd69388: data = 8'he4;
      17'd69389: data = 8'he7;
      17'd69390: data = 8'he5;
      17'd69391: data = 8'hec;
      17'd69392: data = 8'he7;
      17'd69393: data = 8'heb;
      17'd69394: data = 8'h01;
      17'd69395: data = 8'h0e;
      17'd69396: data = 8'h12;
      17'd69397: data = 8'h0e;
      17'd69398: data = 8'h04;
      17'd69399: data = 8'h05;
      17'd69400: data = 8'h0e;
      17'd69401: data = 8'h15;
      17'd69402: data = 8'h19;
      17'd69403: data = 8'h19;
      17'd69404: data = 8'h16;
      17'd69405: data = 8'h11;
      17'd69406: data = 8'h11;
      17'd69407: data = 8'h19;
      17'd69408: data = 8'h16;
      17'd69409: data = 8'h1f;
      17'd69410: data = 8'h27;
      17'd69411: data = 8'h1b;
      17'd69412: data = 8'h1a;
      17'd69413: data = 8'h12;
      17'd69414: data = 8'h13;
      17'd69415: data = 8'h1a;
      17'd69416: data = 8'h16;
      17'd69417: data = 8'h15;
      17'd69418: data = 8'h00;
      17'd69419: data = 8'hf9;
      17'd69420: data = 8'hfa;
      17'd69421: data = 8'hf5;
      17'd69422: data = 8'hfa;
      17'd69423: data = 8'hfe;
      17'd69424: data = 8'hfd;
      17'd69425: data = 8'hfc;
      17'd69426: data = 8'hf4;
      17'd69427: data = 8'hf4;
      17'd69428: data = 8'hf6;
      17'd69429: data = 8'hf6;
      17'd69430: data = 8'hf9;
      17'd69431: data = 8'hf4;
      17'd69432: data = 8'hec;
      17'd69433: data = 8'hec;
      17'd69434: data = 8'hef;
      17'd69435: data = 8'hec;
      17'd69436: data = 8'heb;
      17'd69437: data = 8'he9;
      17'd69438: data = 8'hf1;
      17'd69439: data = 8'hef;
      17'd69440: data = 8'hef;
      17'd69441: data = 8'hfa;
      17'd69442: data = 8'hfd;
      17'd69443: data = 8'h05;
      17'd69444: data = 8'h0c;
      17'd69445: data = 8'h09;
      17'd69446: data = 8'h06;
      17'd69447: data = 8'h05;
      17'd69448: data = 8'h09;
      17'd69449: data = 8'h0d;
      17'd69450: data = 8'h05;
      17'd69451: data = 8'h06;
      17'd69452: data = 8'h09;
      17'd69453: data = 8'h05;
      17'd69454: data = 8'h0a;
      17'd69455: data = 8'h0a;
      17'd69456: data = 8'h0c;
      17'd69457: data = 8'h0e;
      17'd69458: data = 8'h13;
      17'd69459: data = 8'h1b;
      17'd69460: data = 8'h19;
      17'd69461: data = 8'h16;
      17'd69462: data = 8'h16;
      17'd69463: data = 8'h0e;
      17'd69464: data = 8'h0c;
      17'd69465: data = 8'h0a;
      17'd69466: data = 8'h05;
      17'd69467: data = 8'h00;
      17'd69468: data = 8'hfe;
      17'd69469: data = 8'hfe;
      17'd69470: data = 8'hfc;
      17'd69471: data = 8'hf9;
      17'd69472: data = 8'hfa;
      17'd69473: data = 8'hfd;
      17'd69474: data = 8'hfd;
      17'd69475: data = 8'h04;
      17'd69476: data = 8'h04;
      17'd69477: data = 8'h05;
      17'd69478: data = 8'h0c;
      17'd69479: data = 8'h0d;
      17'd69480: data = 8'h06;
      17'd69481: data = 8'h05;
      17'd69482: data = 8'hfe;
      17'd69483: data = 8'hfc;
      17'd69484: data = 8'hfd;
      17'd69485: data = 8'hfe;
      17'd69486: data = 8'hfe;
      17'd69487: data = 8'h0a;
      17'd69488: data = 8'h0e;
      17'd69489: data = 8'h09;
      17'd69490: data = 8'h16;
      17'd69491: data = 8'h16;
      17'd69492: data = 8'h1a;
      17'd69493: data = 8'h27;
      17'd69494: data = 8'h1b;
      17'd69495: data = 8'h1b;
      17'd69496: data = 8'h1f;
      17'd69497: data = 8'h0d;
      17'd69498: data = 8'h11;
      17'd69499: data = 8'h04;
      17'd69500: data = 8'h09;
      17'd69501: data = 8'hfe;
      17'd69502: data = 8'hfa;
      17'd69503: data = 8'h0d;
      17'd69504: data = 8'hfe;
      17'd69505: data = 8'h09;
      17'd69506: data = 8'h0c;
      17'd69507: data = 8'h04;
      17'd69508: data = 8'h0a;
      17'd69509: data = 8'h01;
      17'd69510: data = 8'hf9;
      17'd69511: data = 8'hfd;
      17'd69512: data = 8'hf9;
      17'd69513: data = 8'hfc;
      17'd69514: data = 8'hef;
      17'd69515: data = 8'hec;
      17'd69516: data = 8'he0;
      17'd69517: data = 8'hd6;
      17'd69518: data = 8'he5;
      17'd69519: data = 8'he9;
      17'd69520: data = 8'hf5;
      17'd69521: data = 8'h05;
      17'd69522: data = 8'h05;
      17'd69523: data = 8'h0e;
      17'd69524: data = 8'h12;
      17'd69525: data = 8'h11;
      17'd69526: data = 8'h1a;
      17'd69527: data = 8'h19;
      17'd69528: data = 8'h1b;
      17'd69529: data = 8'h1a;
      17'd69530: data = 8'h13;
      17'd69531: data = 8'h0e;
      17'd69532: data = 8'h01;
      17'd69533: data = 8'h04;
      17'd69534: data = 8'hfe;
      17'd69535: data = 8'hfe;
      17'd69536: data = 8'h01;
      17'd69537: data = 8'hfa;
      17'd69538: data = 8'hf9;
      17'd69539: data = 8'hfe;
      17'd69540: data = 8'h01;
      17'd69541: data = 8'h02;
      17'd69542: data = 8'h0a;
      17'd69543: data = 8'hfd;
      17'd69544: data = 8'hf2;
      17'd69545: data = 8'he4;
      17'd69546: data = 8'hd6;
      17'd69547: data = 8'hd2;
      17'd69548: data = 8'hcb;
      17'd69549: data = 8'hc9;
      17'd69550: data = 8'hc6;
      17'd69551: data = 8'hc5;
      17'd69552: data = 8'hc4;
      17'd69553: data = 8'hbd;
      17'd69554: data = 8'hc0;
      17'd69555: data = 8'hc4;
      17'd69556: data = 8'hca;
      17'd69557: data = 8'hda;
      17'd69558: data = 8'he0;
      17'd69559: data = 8'he2;
      17'd69560: data = 8'he0;
      17'd69561: data = 8'he0;
      17'd69562: data = 8'he0;
      17'd69563: data = 8'he4;
      17'd69564: data = 8'heb;
      17'd69565: data = 8'heb;
      17'd69566: data = 8'hed;
      17'd69567: data = 8'hef;
      17'd69568: data = 8'hf5;
      17'd69569: data = 8'h00;
      17'd69570: data = 8'h0a;
      17'd69571: data = 8'h12;
      17'd69572: data = 8'h1f;
      17'd69573: data = 8'h26;
      17'd69574: data = 8'h29;
      17'd69575: data = 8'h2d;
      17'd69576: data = 8'h31;
      17'd69577: data = 8'h34;
      17'd69578: data = 8'h33;
      17'd69579: data = 8'h33;
      17'd69580: data = 8'h2b;
      17'd69581: data = 8'h22;
      17'd69582: data = 8'h1b;
      17'd69583: data = 8'h12;
      17'd69584: data = 8'h0e;
      17'd69585: data = 8'h11;
      17'd69586: data = 8'h11;
      17'd69587: data = 8'h0e;
      17'd69588: data = 8'h0c;
      17'd69589: data = 8'h04;
      17'd69590: data = 8'h05;
      17'd69591: data = 8'h00;
      17'd69592: data = 8'hfc;
      17'd69593: data = 8'hfa;
      17'd69594: data = 8'hf2;
      17'd69595: data = 8'hed;
      17'd69596: data = 8'he7;
      17'd69597: data = 8'he2;
      17'd69598: data = 8'he0;
      17'd69599: data = 8'hd8;
      17'd69600: data = 8'hd6;
      17'd69601: data = 8'hd6;
      17'd69602: data = 8'hd2;
      17'd69603: data = 8'hd8;
      17'd69604: data = 8'hda;
      17'd69605: data = 8'hde;
      17'd69606: data = 8'he9;
      17'd69607: data = 8'hed;
      17'd69608: data = 8'hf9;
      17'd69609: data = 8'hfe;
      17'd69610: data = 8'hfe;
      17'd69611: data = 8'h02;
      17'd69612: data = 8'h02;
      17'd69613: data = 8'h06;
      17'd69614: data = 8'h0c;
      17'd69615: data = 8'h0d;
      17'd69616: data = 8'h12;
      17'd69617: data = 8'h13;
      17'd69618: data = 8'h13;
      17'd69619: data = 8'h16;
      17'd69620: data = 8'h19;
      17'd69621: data = 8'h1c;
      17'd69622: data = 8'h1f;
      17'd69623: data = 8'h23;
      17'd69624: data = 8'h23;
      17'd69625: data = 8'h23;
      17'd69626: data = 8'h23;
      17'd69627: data = 8'h1f;
      17'd69628: data = 8'h1e;
      17'd69629: data = 8'h19;
      17'd69630: data = 8'h13;
      17'd69631: data = 8'h0d;
      17'd69632: data = 8'h02;
      17'd69633: data = 8'hfd;
      17'd69634: data = 8'hf9;
      17'd69635: data = 8'hf2;
      17'd69636: data = 8'hef;
      17'd69637: data = 8'heb;
      17'd69638: data = 8'he5;
      17'd69639: data = 8'he3;
      17'd69640: data = 8'he2;
      17'd69641: data = 8'he2;
      17'd69642: data = 8'hde;
      17'd69643: data = 8'he0;
      17'd69644: data = 8'he2;
      17'd69645: data = 8'he0;
      17'd69646: data = 8'he2;
      17'd69647: data = 8'he0;
      17'd69648: data = 8'hde;
      17'd69649: data = 8'he0;
      17'd69650: data = 8'he0;
      17'd69651: data = 8'he3;
      17'd69652: data = 8'he4;
      17'd69653: data = 8'he7;
      17'd69654: data = 8'hef;
      17'd69655: data = 8'hf5;
      17'd69656: data = 8'hfe;
      17'd69657: data = 8'h05;
      17'd69658: data = 8'h0c;
      17'd69659: data = 8'h0a;
      17'd69660: data = 8'h09;
      17'd69661: data = 8'h0e;
      17'd69662: data = 8'h0e;
      17'd69663: data = 8'h15;
      17'd69664: data = 8'h23;
      17'd69665: data = 8'h1f;
      17'd69666: data = 8'h1c;
      17'd69667: data = 8'h19;
      17'd69668: data = 8'h0e;
      17'd69669: data = 8'h12;
      17'd69670: data = 8'h12;
      17'd69671: data = 8'h13;
      17'd69672: data = 8'h11;
      17'd69673: data = 8'h0a;
      17'd69674: data = 8'h09;
      17'd69675: data = 8'h09;
      17'd69676: data = 8'h05;
      17'd69677: data = 8'h06;
      17'd69678: data = 8'h05;
      17'd69679: data = 8'h00;
      17'd69680: data = 8'hfa;
      17'd69681: data = 8'hf6;
      17'd69682: data = 8'hf6;
      17'd69683: data = 8'hf9;
      17'd69684: data = 8'hf6;
      17'd69685: data = 8'hf2;
      17'd69686: data = 8'hed;
      17'd69687: data = 8'he2;
      17'd69688: data = 8'he2;
      17'd69689: data = 8'he4;
      17'd69690: data = 8'hec;
      17'd69691: data = 8'hf9;
      17'd69692: data = 8'hfc;
      17'd69693: data = 8'hfd;
      17'd69694: data = 8'h00;
      17'd69695: data = 8'h01;
      17'd69696: data = 8'h05;
      17'd69697: data = 8'h02;
      17'd69698: data = 8'h04;
      17'd69699: data = 8'h05;
      17'd69700: data = 8'h02;
      17'd69701: data = 8'h05;
      17'd69702: data = 8'h02;
      17'd69703: data = 8'h01;
      17'd69704: data = 8'h01;
      17'd69705: data = 8'hfe;
      17'd69706: data = 8'hfe;
      17'd69707: data = 8'hfd;
      17'd69708: data = 8'h00;
      17'd69709: data = 8'h0a;
      17'd69710: data = 8'h0c;
      17'd69711: data = 8'h0e;
      17'd69712: data = 8'h11;
      17'd69713: data = 8'h0e;
      17'd69714: data = 8'h0c;
      17'd69715: data = 8'h05;
      17'd69716: data = 8'h02;
      17'd69717: data = 8'hfe;
      17'd69718: data = 8'hfa;
      17'd69719: data = 8'hfc;
      17'd69720: data = 8'hf6;
      17'd69721: data = 8'hfd;
      17'd69722: data = 8'hfd;
      17'd69723: data = 8'hfc;
      17'd69724: data = 8'h01;
      17'd69725: data = 8'h01;
      17'd69726: data = 8'h05;
      17'd69727: data = 8'h0a;
      17'd69728: data = 8'h0d;
      17'd69729: data = 8'h15;
      17'd69730: data = 8'h12;
      17'd69731: data = 8'h12;
      17'd69732: data = 8'h0d;
      17'd69733: data = 8'h04;
      17'd69734: data = 8'h0a;
      17'd69735: data = 8'h05;
      17'd69736: data = 8'h01;
      17'd69737: data = 8'h0c;
      17'd69738: data = 8'h05;
      17'd69739: data = 8'h05;
      17'd69740: data = 8'h13;
      17'd69741: data = 8'h0a;
      17'd69742: data = 8'h09;
      17'd69743: data = 8'h13;
      17'd69744: data = 8'h0d;
      17'd69745: data = 8'h0d;
      17'd69746: data = 8'h1e;
      17'd69747: data = 8'h13;
      17'd69748: data = 8'h1b;
      17'd69749: data = 8'h29;
      17'd69750: data = 8'h16;
      17'd69751: data = 8'h1c;
      17'd69752: data = 8'h1b;
      17'd69753: data = 8'h0d;
      17'd69754: data = 8'h12;
      17'd69755: data = 8'h19;
      17'd69756: data = 8'h05;
      17'd69757: data = 8'h0e;
      17'd69758: data = 8'h12;
      17'd69759: data = 8'hfd;
      17'd69760: data = 8'h11;
      17'd69761: data = 8'hfe;
      17'd69762: data = 8'hfc;
      17'd69763: data = 8'h19;
      17'd69764: data = 8'hf9;
      17'd69765: data = 8'h04;
      17'd69766: data = 8'h1a;
      17'd69767: data = 8'he9;
      17'd69768: data = 8'h1f;
      17'd69769: data = 8'hfc;
      17'd69770: data = 8'hde;
      17'd69771: data = 8'h16;
      17'd69772: data = 8'hcd;
      17'd69773: data = 8'hf4;
      17'd69774: data = 8'hfa;
      17'd69775: data = 8'hce;
      17'd69776: data = 8'h19;
      17'd69777: data = 8'he5;
      17'd69778: data = 8'h01;
      17'd69779: data = 8'h0d;
      17'd69780: data = 8'he3;
      17'd69781: data = 8'h19;
      17'd69782: data = 8'hf1;
      17'd69783: data = 8'hf9;
      17'd69784: data = 8'h11;
      17'd69785: data = 8'hec;
      17'd69786: data = 8'h11;
      17'd69787: data = 8'h04;
      17'd69788: data = 8'heb;
      17'd69789: data = 8'h0e;
      17'd69790: data = 8'he3;
      17'd69791: data = 8'hfe;
      17'd69792: data = 8'h11;
      17'd69793: data = 8'hfc;
      17'd69794: data = 8'h2d;
      17'd69795: data = 8'h13;
      17'd69796: data = 8'h1a;
      17'd69797: data = 8'h3a;
      17'd69798: data = 8'h02;
      17'd69799: data = 8'h36;
      17'd69800: data = 8'h16;
      17'd69801: data = 8'h11;
      17'd69802: data = 8'h33;
      17'd69803: data = 8'hf5;
      17'd69804: data = 8'h19;
      17'd69805: data = 8'h00;
      17'd69806: data = 8'hec;
      17'd69807: data = 8'h0c;
      17'd69808: data = 8'hd8;
      17'd69809: data = 8'hf4;
      17'd69810: data = 8'heb;
      17'd69811: data = 8'hd2;
      17'd69812: data = 8'hf2;
      17'd69813: data = 8'hdb;
      17'd69814: data = 8'he7;
      17'd69815: data = 8'hf1;
      17'd69816: data = 8'hd5;
      17'd69817: data = 8'he3;
      17'd69818: data = 8'hcd;
      17'd69819: data = 8'hc0;
      17'd69820: data = 8'hce;
      17'd69821: data = 8'hb8;
      17'd69822: data = 8'hc6;
      17'd69823: data = 8'hc6;
      17'd69824: data = 8'hbb;
      17'd69825: data = 8'hcd;
      17'd69826: data = 8'hc0;
      17'd69827: data = 8'hcd;
      17'd69828: data = 8'hd5;
      17'd69829: data = 8'hce;
      17'd69830: data = 8'he9;
      17'd69831: data = 8'he5;
      17'd69832: data = 8'hf6;
      17'd69833: data = 8'hfd;
      17'd69834: data = 8'hf6;
      17'd69835: data = 8'h00;
      17'd69836: data = 8'hfd;
      17'd69837: data = 8'h00;
      17'd69838: data = 8'h02;
      17'd69839: data = 8'h04;
      17'd69840: data = 8'h09;
      17'd69841: data = 8'h0c;
      17'd69842: data = 8'h11;
      17'd69843: data = 8'h16;
      17'd69844: data = 8'h1b;
      17'd69845: data = 8'h1f;
      17'd69846: data = 8'h24;
      17'd69847: data = 8'h22;
      17'd69848: data = 8'h24;
      17'd69849: data = 8'h22;
      17'd69850: data = 8'h1f;
      17'd69851: data = 8'h1f;
      17'd69852: data = 8'h1a;
      17'd69853: data = 8'h1c;
      17'd69854: data = 8'h11;
      17'd69855: data = 8'h0c;
      17'd69856: data = 8'h04;
      17'd69857: data = 8'hf9;
      17'd69858: data = 8'hfc;
      17'd69859: data = 8'hf1;
      17'd69860: data = 8'hf5;
      17'd69861: data = 8'hf6;
      17'd69862: data = 8'hec;
      17'd69863: data = 8'hf6;
      17'd69864: data = 8'heb;
      17'd69865: data = 8'hed;
      17'd69866: data = 8'hef;
      17'd69867: data = 8'he3;
      17'd69868: data = 8'hef;
      17'd69869: data = 8'he3;
      17'd69870: data = 8'he7;
      17'd69871: data = 8'heb;
      17'd69872: data = 8'he3;
      17'd69873: data = 8'hec;
      17'd69874: data = 8'he7;
      17'd69875: data = 8'he9;
      17'd69876: data = 8'hef;
      17'd69877: data = 8'hec;
      17'd69878: data = 8'hf5;
      17'd69879: data = 8'hfa;
      17'd69880: data = 8'h00;
      17'd69881: data = 8'h0c;
      17'd69882: data = 8'h0c;
      17'd69883: data = 8'h11;
      17'd69884: data = 8'h16;
      17'd69885: data = 8'h13;
      17'd69886: data = 8'h1c;
      17'd69887: data = 8'h1b;
      17'd69888: data = 8'h19;
      17'd69889: data = 8'h1e;
      17'd69890: data = 8'h1a;
      17'd69891: data = 8'h1c;
      17'd69892: data = 8'h19;
      17'd69893: data = 8'h12;
      17'd69894: data = 8'h12;
      17'd69895: data = 8'h0a;
      17'd69896: data = 8'h0c;
      17'd69897: data = 8'h0c;
      17'd69898: data = 8'h06;
      17'd69899: data = 8'h09;
      17'd69900: data = 8'h05;
      17'd69901: data = 8'h01;
      17'd69902: data = 8'h00;
      17'd69903: data = 8'hfc;
      17'd69904: data = 8'hf5;
      17'd69905: data = 8'hef;
      17'd69906: data = 8'he9;
      17'd69907: data = 8'he7;
      17'd69908: data = 8'he2;
      17'd69909: data = 8'he0;
      17'd69910: data = 8'hde;
      17'd69911: data = 8'hdb;
      17'd69912: data = 8'hdc;
      17'd69913: data = 8'hdb;
      17'd69914: data = 8'he0;
      17'd69915: data = 8'he2;
      17'd69916: data = 8'he9;
      17'd69917: data = 8'hed;
      17'd69918: data = 8'hef;
      17'd69919: data = 8'hf5;
      17'd69920: data = 8'hf6;
      17'd69921: data = 8'hf9;
      17'd69922: data = 8'hf9;
      17'd69923: data = 8'hfa;
      17'd69924: data = 8'hfd;
      17'd69925: data = 8'hfe;
      17'd69926: data = 8'h01;
      17'd69927: data = 8'h01;
      17'd69928: data = 8'h05;
      17'd69929: data = 8'h06;
      17'd69930: data = 8'h0a;
      17'd69931: data = 8'h0e;
      17'd69932: data = 8'h0e;
      17'd69933: data = 8'h19;
      17'd69934: data = 8'h1a;
      17'd69935: data = 8'h11;
      17'd69936: data = 8'h0d;
      17'd69937: data = 8'h0a;
      17'd69938: data = 8'h05;
      17'd69939: data = 8'h09;
      17'd69940: data = 8'h0d;
      17'd69941: data = 8'h06;
      17'd69942: data = 8'h04;
      17'd69943: data = 8'hfd;
      17'd69944: data = 8'hf4;
      17'd69945: data = 8'hf2;
      17'd69946: data = 8'hf2;
      17'd69947: data = 8'hfa;
      17'd69948: data = 8'hfa;
      17'd69949: data = 8'hf6;
      17'd69950: data = 8'hf2;
      17'd69951: data = 8'he9;
      17'd69952: data = 8'hec;
      17'd69953: data = 8'hf2;
      17'd69954: data = 8'hec;
      17'd69955: data = 8'hed;
      17'd69956: data = 8'hf1;
      17'd69957: data = 8'heb;
      17'd69958: data = 8'hf2;
      17'd69959: data = 8'hfc;
      17'd69960: data = 8'hf9;
      17'd69961: data = 8'hfe;
      17'd69962: data = 8'hfe;
      17'd69963: data = 8'hfa;
      17'd69964: data = 8'hfd;
      17'd69965: data = 8'h01;
      17'd69966: data = 8'h0a;
      17'd69967: data = 8'h11;
      17'd69968: data = 8'h12;
      17'd69969: data = 8'h13;
      17'd69970: data = 8'h0e;
      17'd69971: data = 8'h0c;
      17'd69972: data = 8'h0e;
      17'd69973: data = 8'h0e;
      17'd69974: data = 8'h0d;
      17'd69975: data = 8'h0d;
      17'd69976: data = 8'h0a;
      17'd69977: data = 8'h0a;
      17'd69978: data = 8'h09;
      17'd69979: data = 8'h05;
      17'd69980: data = 8'h05;
      17'd69981: data = 8'h04;
      17'd69982: data = 8'hfe;
      17'd69983: data = 8'hfe;
      17'd69984: data = 8'h00;
      17'd69985: data = 8'hfe;
      17'd69986: data = 8'h01;
      17'd69987: data = 8'h02;
      17'd69988: data = 8'hfe;
      17'd69989: data = 8'hfa;
      17'd69990: data = 8'hf6;
      17'd69991: data = 8'hf4;
      17'd69992: data = 8'hf4;
      17'd69993: data = 8'hfa;
      17'd69994: data = 8'hf9;
      17'd69995: data = 8'hfc;
      17'd69996: data = 8'h01;
      17'd69997: data = 8'h01;
      17'd69998: data = 8'h04;
      17'd69999: data = 8'h04;
      17'd70000: data = 8'h05;
      17'd70001: data = 8'h09;
      17'd70002: data = 8'h09;
      17'd70003: data = 8'h0c;
      17'd70004: data = 8'h0e;
      17'd70005: data = 8'h0e;
      17'd70006: data = 8'h16;
      17'd70007: data = 8'h12;
      17'd70008: data = 8'h0d;
      17'd70009: data = 8'h12;
      17'd70010: data = 8'h0a;
      17'd70011: data = 8'h0c;
      17'd70012: data = 8'h16;
      17'd70013: data = 8'h13;
      17'd70014: data = 8'h0c;
      17'd70015: data = 8'h0c;
      17'd70016: data = 8'h0e;
      17'd70017: data = 8'h09;
      17'd70018: data = 8'h04;
      17'd70019: data = 8'h12;
      17'd70020: data = 8'h04;
      17'd70021: data = 8'h02;
      17'd70022: data = 8'h1b;
      17'd70023: data = 8'h01;
      17'd70024: data = 8'h04;
      17'd70025: data = 8'h19;
      17'd70026: data = 8'h02;
      17'd70027: data = 8'h0c;
      17'd70028: data = 8'h05;
      17'd70029: data = 8'h01;
      17'd70030: data = 8'h00;
      17'd70031: data = 8'hf6;
      17'd70032: data = 8'h01;
      17'd70033: data = 8'hed;
      17'd70034: data = 8'hf9;
      17'd70035: data = 8'h02;
      17'd70036: data = 8'hf9;
      17'd70037: data = 8'h11;
      17'd70038: data = 8'h01;
      17'd70039: data = 8'h0c;
      17'd70040: data = 8'h1e;
      17'd70041: data = 8'h04;
      17'd70042: data = 8'h11;
      17'd70043: data = 8'h0d;
      17'd70044: data = 8'h05;
      17'd70045: data = 8'h0d;
      17'd70046: data = 8'hfd;
      17'd70047: data = 8'h0c;
      17'd70048: data = 8'hf4;
      17'd70049: data = 8'hf5;
      17'd70050: data = 8'h0e;
      17'd70051: data = 8'hf6;
      17'd70052: data = 8'hfe;
      17'd70053: data = 8'h0d;
      17'd70054: data = 8'h06;
      17'd70055: data = 8'h09;
      17'd70056: data = 8'h0d;
      17'd70057: data = 8'h0d;
      17'd70058: data = 8'h04;
      17'd70059: data = 8'hfc;
      17'd70060: data = 8'h00;
      17'd70061: data = 8'h00;
      17'd70062: data = 8'hed;
      17'd70063: data = 8'h02;
      17'd70064: data = 8'hfe;
      17'd70065: data = 8'hef;
      17'd70066: data = 8'hfd;
      17'd70067: data = 8'hde;
      17'd70068: data = 8'hfa;
      17'd70069: data = 8'hf1;
      17'd70070: data = 8'hed;
      17'd70071: data = 8'h0a;
      17'd70072: data = 8'hf2;
      17'd70073: data = 8'h0c;
      17'd70074: data = 8'h05;
      17'd70075: data = 8'h02;
      17'd70076: data = 8'h12;
      17'd70077: data = 8'hfc;
      17'd70078: data = 8'h13;
      17'd70079: data = 8'h04;
      17'd70080: data = 8'hf6;
      17'd70081: data = 8'h04;
      17'd70082: data = 8'hfd;
      17'd70083: data = 8'hfe;
      17'd70084: data = 8'h06;
      17'd70085: data = 8'hfe;
      17'd70086: data = 8'hf9;
      17'd70087: data = 8'hf4;
      17'd70088: data = 8'hed;
      17'd70089: data = 8'hfc;
      17'd70090: data = 8'hfa;
      17'd70091: data = 8'h00;
      17'd70092: data = 8'h00;
      17'd70093: data = 8'hf1;
      17'd70094: data = 8'hfc;
      17'd70095: data = 8'hec;
      17'd70096: data = 8'he7;
      17'd70097: data = 8'hf1;
      17'd70098: data = 8'hda;
      17'd70099: data = 8'he4;
      17'd70100: data = 8'hdb;
      17'd70101: data = 8'hda;
      17'd70102: data = 8'he3;
      17'd70103: data = 8'hd6;
      17'd70104: data = 8'hde;
      17'd70105: data = 8'hdc;
      17'd70106: data = 8'hdb;
      17'd70107: data = 8'he2;
      17'd70108: data = 8'hde;
      17'd70109: data = 8'he5;
      17'd70110: data = 8'hed;
      17'd70111: data = 8'hec;
      17'd70112: data = 8'hf4;
      17'd70113: data = 8'hf1;
      17'd70114: data = 8'hec;
      17'd70115: data = 8'hf5;
      17'd70116: data = 8'hf1;
      17'd70117: data = 8'hf6;
      17'd70118: data = 8'hf9;
      17'd70119: data = 8'hf9;
      17'd70120: data = 8'h04;
      17'd70121: data = 8'hfe;
      17'd70122: data = 8'h0c;
      17'd70123: data = 8'h0d;
      17'd70124: data = 8'h0a;
      17'd70125: data = 8'h12;
      17'd70126: data = 8'h0d;
      17'd70127: data = 8'h13;
      17'd70128: data = 8'h19;
      17'd70129: data = 8'h1e;
      17'd70130: data = 8'h23;
      17'd70131: data = 8'h1b;
      17'd70132: data = 8'h1a;
      17'd70133: data = 8'h12;
      17'd70134: data = 8'h11;
      17'd70135: data = 8'h0e;
      17'd70136: data = 8'h0c;
      17'd70137: data = 8'h06;
      17'd70138: data = 8'h06;
      17'd70139: data = 8'h04;
      17'd70140: data = 8'h01;
      17'd70141: data = 8'h06;
      17'd70142: data = 8'h02;
      17'd70143: data = 8'h02;
      17'd70144: data = 8'h00;
      17'd70145: data = 8'hfd;
      17'd70146: data = 8'hfe;
      17'd70147: data = 8'hfa;
      17'd70148: data = 8'hfe;
      17'd70149: data = 8'hfc;
      17'd70150: data = 8'hf9;
      17'd70151: data = 8'hf6;
      17'd70152: data = 8'hef;
      17'd70153: data = 8'hef;
      17'd70154: data = 8'he9;
      17'd70155: data = 8'hef;
      17'd70156: data = 8'hf4;
      17'd70157: data = 8'hf4;
      17'd70158: data = 8'hf9;
      17'd70159: data = 8'hfa;
      17'd70160: data = 8'h00;
      17'd70161: data = 8'h02;
      17'd70162: data = 8'h04;
      17'd70163: data = 8'h06;
      17'd70164: data = 8'h09;
      17'd70165: data = 8'h09;
      17'd70166: data = 8'h0c;
      17'd70167: data = 8'h0c;
      17'd70168: data = 8'h0c;
      17'd70169: data = 8'h0e;
      17'd70170: data = 8'h0a;
      17'd70171: data = 8'h09;
      17'd70172: data = 8'h05;
      17'd70173: data = 8'h05;
      17'd70174: data = 8'h0c;
      17'd70175: data = 8'h0c;
      17'd70176: data = 8'h0d;
      17'd70177: data = 8'h0c;
      17'd70178: data = 8'h0d;
      17'd70179: data = 8'h0d;
      17'd70180: data = 8'h06;
      17'd70181: data = 8'h0a;
      17'd70182: data = 8'h04;
      17'd70183: data = 8'h01;
      17'd70184: data = 8'h01;
      17'd70185: data = 8'hfd;
      17'd70186: data = 8'hfc;
      17'd70187: data = 8'hfa;
      17'd70188: data = 8'hf5;
      17'd70189: data = 8'hf4;
      17'd70190: data = 8'hef;
      17'd70191: data = 8'hef;
      17'd70192: data = 8'hef;
      17'd70193: data = 8'hf1;
      17'd70194: data = 8'hf2;
      17'd70195: data = 8'hf2;
      17'd70196: data = 8'hf2;
      17'd70197: data = 8'hf4;
      17'd70198: data = 8'hf2;
      17'd70199: data = 8'hf4;
      17'd70200: data = 8'hf4;
      17'd70201: data = 8'hf2;
      17'd70202: data = 8'hf5;
      17'd70203: data = 8'hf4;
      17'd70204: data = 8'hf5;
      17'd70205: data = 8'hf6;
      17'd70206: data = 8'hf9;
      17'd70207: data = 8'hfc;
      17'd70208: data = 8'hfc;
      17'd70209: data = 8'hfe;
      17'd70210: data = 8'hfd;
      17'd70211: data = 8'hfe;
      17'd70212: data = 8'h04;
      17'd70213: data = 8'h06;
      17'd70214: data = 8'h0d;
      17'd70215: data = 8'h0c;
      17'd70216: data = 8'h00;
      17'd70217: data = 8'hfe;
      17'd70218: data = 8'hfa;
      17'd70219: data = 8'hf6;
      17'd70220: data = 8'h05;
      17'd70221: data = 8'h0c;
      17'd70222: data = 8'h06;
      17'd70223: data = 8'h09;
      17'd70224: data = 8'h02;
      17'd70225: data = 8'hfc;
      17'd70226: data = 8'h01;
      17'd70227: data = 8'h05;
      17'd70228: data = 8'h05;
      17'd70229: data = 8'h01;
      17'd70230: data = 8'hfe;
      17'd70231: data = 8'hf9;
      17'd70232: data = 8'hf5;
      17'd70233: data = 8'hfd;
      17'd70234: data = 8'hfd;
      17'd70235: data = 8'hf9;
      17'd70236: data = 8'hfd;
      17'd70237: data = 8'hf9;
      17'd70238: data = 8'hf2;
      17'd70239: data = 8'hfa;
      17'd70240: data = 8'hfe;
      17'd70241: data = 8'h01;
      17'd70242: data = 8'h04;
      17'd70243: data = 8'h04;
      17'd70244: data = 8'hfe;
      17'd70245: data = 8'hfe;
      17'd70246: data = 8'h06;
      17'd70247: data = 8'h09;
      17'd70248: data = 8'h09;
      17'd70249: data = 8'h0d;
      17'd70250: data = 8'h05;
      17'd70251: data = 8'h04;
      17'd70252: data = 8'h05;
      17'd70253: data = 8'h04;
      17'd70254: data = 8'h05;
      17'd70255: data = 8'h02;
      17'd70256: data = 8'h00;
      17'd70257: data = 8'h00;
      17'd70258: data = 8'hfd;
      17'd70259: data = 8'hfe;
      17'd70260: data = 8'hfe;
      17'd70261: data = 8'h02;
      17'd70262: data = 8'h04;
      17'd70263: data = 8'hfe;
      17'd70264: data = 8'hfd;
      17'd70265: data = 8'hfe;
      17'd70266: data = 8'hfd;
      17'd70267: data = 8'h00;
      17'd70268: data = 8'h00;
      17'd70269: data = 8'hfe;
      17'd70270: data = 8'hfc;
      17'd70271: data = 8'hf6;
      17'd70272: data = 8'hfa;
      17'd70273: data = 8'hfc;
      17'd70274: data = 8'h00;
      17'd70275: data = 8'h01;
      17'd70276: data = 8'h01;
      17'd70277: data = 8'h00;
      17'd70278: data = 8'h01;
      17'd70279: data = 8'h06;
      17'd70280: data = 8'h0c;
      17'd70281: data = 8'h09;
      17'd70282: data = 8'h0c;
      17'd70283: data = 8'h0c;
      17'd70284: data = 8'h06;
      17'd70285: data = 8'h0d;
      17'd70286: data = 8'h0e;
      17'd70287: data = 8'h11;
      17'd70288: data = 8'h0d;
      17'd70289: data = 8'h0a;
      17'd70290: data = 8'h06;
      17'd70291: data = 8'h06;
      17'd70292: data = 8'h09;
      17'd70293: data = 8'h0d;
      17'd70294: data = 8'h0d;
      17'd70295: data = 8'h0c;
      17'd70296: data = 8'h0c;
      17'd70297: data = 8'h0a;
      17'd70298: data = 8'h06;
      17'd70299: data = 8'h05;
      17'd70300: data = 8'h0a;
      17'd70301: data = 8'h00;
      17'd70302: data = 8'hfe;
      17'd70303: data = 8'h05;
      17'd70304: data = 8'h04;
      17'd70305: data = 8'h0a;
      17'd70306: data = 8'h13;
      17'd70307: data = 8'h0d;
      17'd70308: data = 8'h12;
      17'd70309: data = 8'h05;
      17'd70310: data = 8'h00;
      17'd70311: data = 8'h13;
      17'd70312: data = 8'hfc;
      17'd70313: data = 8'hfa;
      17'd70314: data = 8'h13;
      17'd70315: data = 8'hf4;
      17'd70316: data = 8'hf2;
      17'd70317: data = 8'h23;
      17'd70318: data = 8'hf1;
      17'd70319: data = 8'h00;
      17'd70320: data = 8'h23;
      17'd70321: data = 8'heb;
      17'd70322: data = 8'h0c;
      17'd70323: data = 8'h09;
      17'd70324: data = 8'hf5;
      17'd70325: data = 8'h1a;
      17'd70326: data = 8'hf4;
      17'd70327: data = 8'h06;
      17'd70328: data = 8'h0e;
      17'd70329: data = 8'hd8;
      17'd70330: data = 8'h11;
      17'd70331: data = 8'hf6;
      17'd70332: data = 8'hf4;
      17'd70333: data = 8'h06;
      17'd70334: data = 8'hf6;
      17'd70335: data = 8'h04;
      17'd70336: data = 8'hfa;
      17'd70337: data = 8'h05;
      17'd70338: data = 8'h02;
      17'd70339: data = 8'he7;
      17'd70340: data = 8'hf5;
      17'd70341: data = 8'he4;
      17'd70342: data = 8'hdb;
      17'd70343: data = 8'hf9;
      17'd70344: data = 8'h01;
      17'd70345: data = 8'h01;
      17'd70346: data = 8'h13;
      17'd70347: data = 8'h16;
      17'd70348: data = 8'hfe;
      17'd70349: data = 8'h0c;
      17'd70350: data = 8'h13;
      17'd70351: data = 8'h12;
      17'd70352: data = 8'h06;
      17'd70353: data = 8'h05;
      17'd70354: data = 8'h16;
      17'd70355: data = 8'he9;
      17'd70356: data = 8'h0d;
      17'd70357: data = 8'h02;
      17'd70358: data = 8'heb;
      17'd70359: data = 8'h12;
      17'd70360: data = 8'he7;
      17'd70361: data = 8'h00;
      17'd70362: data = 8'hfd;
      17'd70363: data = 8'h04;
      17'd70364: data = 8'h1b;
      17'd70365: data = 8'h04;
      17'd70366: data = 8'h12;
      17'd70367: data = 8'h01;
      17'd70368: data = 8'hef;
      17'd70369: data = 8'h0c;
      17'd70370: data = 8'hf1;
      17'd70371: data = 8'hf4;
      17'd70372: data = 8'hf5;
      17'd70373: data = 8'he4;
      17'd70374: data = 8'he3;
      17'd70375: data = 8'he3;
      17'd70376: data = 8'he4;
      17'd70377: data = 8'he3;
      17'd70378: data = 8'he0;
      17'd70379: data = 8'he3;
      17'd70380: data = 8'he2;
      17'd70381: data = 8'hd8;
      17'd70382: data = 8'hf5;
      17'd70383: data = 8'hed;
      17'd70384: data = 8'hef;
      17'd70385: data = 8'hf5;
      17'd70386: data = 8'hdb;
      17'd70387: data = 8'heb;
      17'd70388: data = 8'he3;
      17'd70389: data = 8'he3;
      17'd70390: data = 8'hf4;
      17'd70391: data = 8'he4;
      17'd70392: data = 8'hf1;
      17'd70393: data = 8'he9;
      17'd70394: data = 8'he0;
      17'd70395: data = 8'hf6;
      17'd70396: data = 8'he9;
      17'd70397: data = 8'hfa;
      17'd70398: data = 8'h02;
      17'd70399: data = 8'hf5;
      17'd70400: data = 8'h0a;
      17'd70401: data = 8'h02;
      17'd70402: data = 8'h0a;
      17'd70403: data = 8'h12;
      17'd70404: data = 8'h06;
      17'd70405: data = 8'h0d;
      17'd70406: data = 8'h04;
      17'd70407: data = 8'h00;
      17'd70408: data = 8'h05;
      17'd70409: data = 8'h01;
      17'd70410: data = 8'h0a;
      17'd70411: data = 8'h06;
      17'd70412: data = 8'hfe;
      17'd70413: data = 8'h05;
      17'd70414: data = 8'h00;
      17'd70415: data = 8'h04;
      17'd70416: data = 8'h0e;
      17'd70417: data = 8'h06;
      17'd70418: data = 8'h0c;
      17'd70419: data = 8'h0c;
      17'd70420: data = 8'h02;
      17'd70421: data = 8'h0d;
      17'd70422: data = 8'h00;
      17'd70423: data = 8'h01;
      17'd70424: data = 8'hfe;
      17'd70425: data = 8'hf2;
      17'd70426: data = 8'hfc;
      17'd70427: data = 8'hed;
      17'd70428: data = 8'hf9;
      17'd70429: data = 8'hfa;
      17'd70430: data = 8'hf1;
      17'd70431: data = 8'hfd;
      17'd70432: data = 8'hf6;
      17'd70433: data = 8'hf6;
      17'd70434: data = 8'hfe;
      17'd70435: data = 8'hfc;
      17'd70436: data = 8'h04;
      17'd70437: data = 8'h04;
      17'd70438: data = 8'h01;
      17'd70439: data = 8'h06;
      17'd70440: data = 8'hfe;
      17'd70441: data = 8'h01;
      17'd70442: data = 8'h04;
      17'd70443: data = 8'hfe;
      17'd70444: data = 8'h01;
      17'd70445: data = 8'hfd;
      17'd70446: data = 8'hfe;
      17'd70447: data = 8'h05;
      17'd70448: data = 8'h02;
      17'd70449: data = 8'h06;
      17'd70450: data = 8'h09;
      17'd70451: data = 8'h04;
      17'd70452: data = 8'h0a;
      17'd70453: data = 8'h09;
      17'd70454: data = 8'h0c;
      17'd70455: data = 8'h0c;
      17'd70456: data = 8'h09;
      17'd70457: data = 8'h0a;
      17'd70458: data = 8'h04;
      17'd70459: data = 8'h00;
      17'd70460: data = 8'h04;
      17'd70461: data = 8'hfc;
      17'd70462: data = 8'hfd;
      17'd70463: data = 8'hfc;
      17'd70464: data = 8'hf4;
      17'd70465: data = 8'hfa;
      17'd70466: data = 8'hf6;
      17'd70467: data = 8'hfc;
      17'd70468: data = 8'hfe;
      17'd70469: data = 8'hfc;
      17'd70470: data = 8'h01;
      17'd70471: data = 8'hfc;
      17'd70472: data = 8'hfe;
      17'd70473: data = 8'h02;
      17'd70474: data = 8'hfa;
      17'd70475: data = 8'hfe;
      17'd70476: data = 8'hfd;
      17'd70477: data = 8'hf5;
      17'd70478: data = 8'hf5;
      17'd70479: data = 8'hf4;
      17'd70480: data = 8'hf4;
      17'd70481: data = 8'hf5;
      17'd70482: data = 8'hf6;
      17'd70483: data = 8'hf9;
      17'd70484: data = 8'hfa;
      17'd70485: data = 8'hfc;
      17'd70486: data = 8'hfe;
      17'd70487: data = 8'hfe;
      17'd70488: data = 8'h01;
      17'd70489: data = 8'h04;
      17'd70490: data = 8'h00;
      17'd70491: data = 8'hfe;
      17'd70492: data = 8'h00;
      17'd70493: data = 8'hfd;
      17'd70494: data = 8'hfe;
      17'd70495: data = 8'h00;
      17'd70496: data = 8'hfc;
      17'd70497: data = 8'hf5;
      17'd70498: data = 8'hf6;
      17'd70499: data = 8'hf9;
      17'd70500: data = 8'hf2;
      17'd70501: data = 8'h01;
      17'd70502: data = 8'h01;
      17'd70503: data = 8'hf2;
      17'd70504: data = 8'hfd;
      17'd70505: data = 8'hfd;
      17'd70506: data = 8'hf6;
      17'd70507: data = 8'h01;
      17'd70508: data = 8'h09;
      17'd70509: data = 8'h01;
      17'd70510: data = 8'hfd;
      17'd70511: data = 8'h00;
      17'd70512: data = 8'h02;
      17'd70513: data = 8'h00;
      17'd70514: data = 8'h05;
      17'd70515: data = 8'h09;
      17'd70516: data = 8'hfa;
      17'd70517: data = 8'hfc;
      17'd70518: data = 8'hfe;
      17'd70519: data = 8'hf6;
      17'd70520: data = 8'h01;
      17'd70521: data = 8'h06;
      17'd70522: data = 8'h00;
      17'd70523: data = 8'hfd;
      17'd70524: data = 8'h02;
      17'd70525: data = 8'h04;
      17'd70526: data = 8'h04;
      17'd70527: data = 8'h0d;
      17'd70528: data = 8'h13;
      17'd70529: data = 8'h04;
      17'd70530: data = 8'h04;
      17'd70531: data = 8'h06;
      17'd70532: data = 8'h02;
      17'd70533: data = 8'h05;
      17'd70534: data = 8'h05;
      17'd70535: data = 8'h01;
      17'd70536: data = 8'h00;
      17'd70537: data = 8'hfc;
      17'd70538: data = 8'hfc;
      17'd70539: data = 8'hfc;
      17'd70540: data = 8'hfd;
      17'd70541: data = 8'h01;
      17'd70542: data = 8'h00;
      17'd70543: data = 8'h00;
      17'd70544: data = 8'hfe;
      17'd70545: data = 8'hfd;
      17'd70546: data = 8'h01;
      17'd70547: data = 8'h01;
      17'd70548: data = 8'hfd;
      17'd70549: data = 8'hfe;
      17'd70550: data = 8'hfd;
      17'd70551: data = 8'hfa;
      17'd70552: data = 8'hfc;
      17'd70553: data = 8'hfe;
      17'd70554: data = 8'hfc;
      17'd70555: data = 8'hfc;
      17'd70556: data = 8'hfd;
      17'd70557: data = 8'hfe;
      17'd70558: data = 8'hfe;
      17'd70559: data = 8'h01;
      17'd70560: data = 8'h05;
      17'd70561: data = 8'h06;
      17'd70562: data = 8'h06;
      17'd70563: data = 8'h04;
      17'd70564: data = 8'h04;
      17'd70565: data = 8'h06;
      17'd70566: data = 8'h0a;
      17'd70567: data = 8'h09;
      17'd70568: data = 8'h09;
      17'd70569: data = 8'h06;
      17'd70570: data = 8'h04;
      17'd70571: data = 8'h09;
      17'd70572: data = 8'h09;
      17'd70573: data = 8'h0c;
      17'd70574: data = 8'h11;
      17'd70575: data = 8'h0a;
      17'd70576: data = 8'h09;
      17'd70577: data = 8'h0a;
      17'd70578: data = 8'h09;
      17'd70579: data = 8'h06;
      17'd70580: data = 8'h06;
      17'd70581: data = 8'h09;
      17'd70582: data = 8'h05;
      17'd70583: data = 8'h01;
      17'd70584: data = 8'h06;
      17'd70585: data = 8'h09;
      17'd70586: data = 8'h04;
      17'd70587: data = 8'h0a;
      17'd70588: data = 8'h0d;
      17'd70589: data = 8'h05;
      17'd70590: data = 8'h06;
      17'd70591: data = 8'h09;
      17'd70592: data = 8'h06;
      17'd70593: data = 8'h05;
      17'd70594: data = 8'h0a;
      17'd70595: data = 8'h0c;
      17'd70596: data = 8'hf9;
      17'd70597: data = 8'h01;
      17'd70598: data = 8'h09;
      17'd70599: data = 8'hef;
      17'd70600: data = 8'h09;
      17'd70601: data = 8'h15;
      17'd70602: data = 8'hec;
      17'd70603: data = 8'h09;
      17'd70604: data = 8'h0e;
      17'd70605: data = 8'hf2;
      17'd70606: data = 8'h0a;
      17'd70607: data = 8'h06;
      17'd70608: data = 8'hfe;
      17'd70609: data = 8'h02;
      17'd70610: data = 8'h00;
      17'd70611: data = 8'h0a;
      17'd70612: data = 8'h09;
      17'd70613: data = 8'h05;
      17'd70614: data = 8'h06;
      17'd70615: data = 8'h05;
      17'd70616: data = 8'hfe;
      17'd70617: data = 8'h06;
      17'd70618: data = 8'h11;
      17'd70619: data = 8'h06;
      17'd70620: data = 8'h09;
      17'd70621: data = 8'hf2;
      17'd70622: data = 8'hf4;
      17'd70623: data = 8'he0;
      17'd70624: data = 8'hec;
      17'd70625: data = 8'hf9;
      17'd70626: data = 8'hf4;
      17'd70627: data = 8'h02;
      17'd70628: data = 8'h01;
      17'd70629: data = 8'h06;
      17'd70630: data = 8'h02;
      17'd70631: data = 8'h0e;
      17'd70632: data = 8'h11;
      17'd70633: data = 8'hfa;
      17'd70634: data = 8'h04;
      17'd70635: data = 8'hf9;
      17'd70636: data = 8'he5;
      17'd70637: data = 8'hf6;
      17'd70638: data = 8'hf2;
      17'd70639: data = 8'heb;
      17'd70640: data = 8'he2;
      17'd70641: data = 8'heb;
      17'd70642: data = 8'heb;
      17'd70643: data = 8'hde;
      17'd70644: data = 8'hfe;
      17'd70645: data = 8'h00;
      17'd70646: data = 8'h04;
      17'd70647: data = 8'h01;
      17'd70648: data = 8'h0c;
      17'd70649: data = 8'hfd;
      17'd70650: data = 8'hfa;
      17'd70651: data = 8'h02;
      17'd70652: data = 8'hf5;
      17'd70653: data = 8'hfc;
      17'd70654: data = 8'hef;
      17'd70655: data = 8'hf9;
      17'd70656: data = 8'heb;
      17'd70657: data = 8'hf4;
      17'd70658: data = 8'hf6;
      17'd70659: data = 8'hec;
      17'd70660: data = 8'hf4;
      17'd70661: data = 8'hf9;
      17'd70662: data = 8'hf5;
      17'd70663: data = 8'h02;
      17'd70664: data = 8'h05;
      17'd70665: data = 8'h09;
      17'd70666: data = 8'h05;
      17'd70667: data = 8'hfd;
      17'd70668: data = 8'h04;
      17'd70669: data = 8'hf2;
      17'd70670: data = 8'hfa;
      17'd70671: data = 8'hf6;
      17'd70672: data = 8'hf5;
      17'd70673: data = 8'hf5;
      17'd70674: data = 8'hef;
      17'd70675: data = 8'hef;
      17'd70676: data = 8'hed;
      17'd70677: data = 8'hf1;
      17'd70678: data = 8'heb;
      17'd70679: data = 8'hf6;
      17'd70680: data = 8'hf1;
      17'd70681: data = 8'hf5;
      17'd70682: data = 8'hf6;
      17'd70683: data = 8'hf9;
      17'd70684: data = 8'hfa;
      17'd70685: data = 8'hf5;
      17'd70686: data = 8'hf6;
      17'd70687: data = 8'hf1;
      17'd70688: data = 8'hf2;
      17'd70689: data = 8'hf5;
      17'd70690: data = 8'hf4;
      17'd70691: data = 8'hf5;
      17'd70692: data = 8'hf9;
      17'd70693: data = 8'hf2;
      17'd70694: data = 8'hf5;
      17'd70695: data = 8'hf6;
      17'd70696: data = 8'hfa;
      17'd70697: data = 8'hfc;
      17'd70698: data = 8'h01;
      17'd70699: data = 8'h04;
      17'd70700: data = 8'h00;
      17'd70701: data = 8'h04;
      17'd70702: data = 8'h06;
      17'd70703: data = 8'h04;
      17'd70704: data = 8'h05;
      17'd70705: data = 8'h06;
      17'd70706: data = 8'h00;
      17'd70707: data = 8'h02;
      17'd70708: data = 8'h02;
      17'd70709: data = 8'hfe;
      17'd70710: data = 8'h01;
      17'd70711: data = 8'h00;
      17'd70712: data = 8'h00;
      17'd70713: data = 8'hfd;
      17'd70714: data = 8'hfe;
      17'd70715: data = 8'h04;
      17'd70716: data = 8'h02;
      17'd70717: data = 8'h0a;
      17'd70718: data = 8'h0d;
      17'd70719: data = 8'h06;
      17'd70720: data = 8'h05;
      17'd70721: data = 8'h04;
      17'd70722: data = 8'h05;
      17'd70723: data = 8'h00;
      17'd70724: data = 8'hfe;
      17'd70725: data = 8'hfe;
      17'd70726: data = 8'hfc;
      17'd70727: data = 8'hfd;
      17'd70728: data = 8'hfd;
      17'd70729: data = 8'hfd;
      17'd70730: data = 8'hfe;
      17'd70731: data = 8'hfe;
      17'd70732: data = 8'hfd;
      17'd70733: data = 8'h01;
      17'd70734: data = 8'h02;
      17'd70735: data = 8'h04;
      17'd70736: data = 8'h04;
      17'd70737: data = 8'h05;
      17'd70738: data = 8'h02;
      17'd70739: data = 8'h00;
      17'd70740: data = 8'hfe;
      17'd70741: data = 8'h00;
      17'd70742: data = 8'h00;
      17'd70743: data = 8'hfe;
      17'd70744: data = 8'hfe;
      17'd70745: data = 8'hfd;
      17'd70746: data = 8'h00;
      17'd70747: data = 8'hfe;
      17'd70748: data = 8'h01;
      17'd70749: data = 8'h02;
      17'd70750: data = 8'h00;
      17'd70751: data = 8'h02;
      17'd70752: data = 8'h02;
      17'd70753: data = 8'h02;
      17'd70754: data = 8'h05;
      17'd70755: data = 8'h06;
      17'd70756: data = 8'h06;
      17'd70757: data = 8'hfe;
      17'd70758: data = 8'hfe;
      17'd70759: data = 8'hfe;
      17'd70760: data = 8'hfd;
      17'd70761: data = 8'h00;
      17'd70762: data = 8'h02;
      17'd70763: data = 8'hfc;
      17'd70764: data = 8'hfc;
      17'd70765: data = 8'hfe;
      17'd70766: data = 8'hfd;
      17'd70767: data = 8'hfd;
      17'd70768: data = 8'hfe;
      17'd70769: data = 8'hfe;
      17'd70770: data = 8'hfc;
      17'd70771: data = 8'hfd;
      17'd70772: data = 8'h01;
      17'd70773: data = 8'h00;
      17'd70774: data = 8'hfe;
      17'd70775: data = 8'h02;
      17'd70776: data = 8'hfd;
      17'd70777: data = 8'hf5;
      17'd70778: data = 8'hf9;
      17'd70779: data = 8'hfa;
      17'd70780: data = 8'hf9;
      17'd70781: data = 8'h00;
      17'd70782: data = 8'h01;
      17'd70783: data = 8'hfd;
      17'd70784: data = 8'hf9;
      17'd70785: data = 8'hf1;
      17'd70786: data = 8'hf6;
      17'd70787: data = 8'hfe;
      17'd70788: data = 8'hf9;
      17'd70789: data = 8'hfd;
      17'd70790: data = 8'h00;
      17'd70791: data = 8'hf5;
      17'd70792: data = 8'hfe;
      17'd70793: data = 8'h06;
      17'd70794: data = 8'h04;
      17'd70795: data = 8'h0e;
      17'd70796: data = 8'h0a;
      17'd70797: data = 8'h04;
      17'd70798: data = 8'h01;
      17'd70799: data = 8'h02;
      17'd70800: data = 8'h09;
      17'd70801: data = 8'h04;
      17'd70802: data = 8'h01;
      17'd70803: data = 8'h04;
      17'd70804: data = 8'hfd;
      17'd70805: data = 8'hf6;
      17'd70806: data = 8'h00;
      17'd70807: data = 8'h04;
      17'd70808: data = 8'hfe;
      17'd70809: data = 8'h02;
      17'd70810: data = 8'h00;
      17'd70811: data = 8'hfc;
      17'd70812: data = 8'h00;
      17'd70813: data = 8'h00;
      17'd70814: data = 8'h02;
      17'd70815: data = 8'hfe;
      17'd70816: data = 8'hfc;
      17'd70817: data = 8'hfc;
      17'd70818: data = 8'hf9;
      17'd70819: data = 8'hfd;
      17'd70820: data = 8'hfe;
      17'd70821: data = 8'hfe;
      17'd70822: data = 8'h02;
      17'd70823: data = 8'hfd;
      17'd70824: data = 8'hfa;
      17'd70825: data = 8'hfd;
      17'd70826: data = 8'hfe;
      17'd70827: data = 8'h01;
      17'd70828: data = 8'h02;
      17'd70829: data = 8'h01;
      17'd70830: data = 8'h01;
      17'd70831: data = 8'h01;
      17'd70832: data = 8'h00;
      17'd70833: data = 8'h02;
      17'd70834: data = 8'h05;
      17'd70835: data = 8'h04;
      17'd70836: data = 8'h01;
      17'd70837: data = 8'h02;
      17'd70838: data = 8'h06;
      17'd70839: data = 8'h04;
      17'd70840: data = 8'h02;
      17'd70841: data = 8'h06;
      17'd70842: data = 8'h05;
      17'd70843: data = 8'h02;
      17'd70844: data = 8'h02;
      17'd70845: data = 8'h06;
      17'd70846: data = 8'h09;
      17'd70847: data = 8'h09;
      17'd70848: data = 8'h0d;
      17'd70849: data = 8'h09;
      17'd70850: data = 8'h05;
      17'd70851: data = 8'h0a;
      17'd70852: data = 8'h0a;
      17'd70853: data = 8'h09;
      17'd70854: data = 8'h0c;
      17'd70855: data = 8'h09;
      17'd70856: data = 8'h04;
      17'd70857: data = 8'h06;
      17'd70858: data = 8'h06;
      17'd70859: data = 8'h05;
      17'd70860: data = 8'h06;
      17'd70861: data = 8'h09;
      17'd70862: data = 8'h06;
      17'd70863: data = 8'h04;
      17'd70864: data = 8'h09;
      17'd70865: data = 8'h0a;
      17'd70866: data = 8'h0a;
      17'd70867: data = 8'h0d;
      17'd70868: data = 8'h09;
      17'd70869: data = 8'h02;
      17'd70870: data = 8'h02;
      17'd70871: data = 8'h04;
      17'd70872: data = 8'h04;
      17'd70873: data = 8'h02;
      17'd70874: data = 8'h04;
      17'd70875: data = 8'h02;
      17'd70876: data = 8'hfe;
      17'd70877: data = 8'h00;
      17'd70878: data = 8'h00;
      17'd70879: data = 8'h00;
      17'd70880: data = 8'h01;
      17'd70881: data = 8'h04;
      17'd70882: data = 8'h04;
      17'd70883: data = 8'h01;
      17'd70884: data = 8'h06;
      17'd70885: data = 8'h04;
      17'd70886: data = 8'h00;
      17'd70887: data = 8'h05;
      17'd70888: data = 8'h02;
      17'd70889: data = 8'hfe;
      17'd70890: data = 8'h04;
      17'd70891: data = 8'h04;
      17'd70892: data = 8'h02;
      17'd70893: data = 8'h02;
      17'd70894: data = 8'h02;
      17'd70895: data = 8'h00;
      17'd70896: data = 8'h00;
      17'd70897: data = 8'h04;
      17'd70898: data = 8'h04;
      17'd70899: data = 8'h02;
      17'd70900: data = 8'h0e;
      17'd70901: data = 8'h0d;
      17'd70902: data = 8'h02;
      17'd70903: data = 8'h11;
      17'd70904: data = 8'h13;
      17'd70905: data = 8'hfd;
      17'd70906: data = 8'h0c;
      17'd70907: data = 8'h09;
      17'd70908: data = 8'hf2;
      17'd70909: data = 8'hfe;
      17'd70910: data = 8'h02;
      17'd70911: data = 8'hf5;
      17'd70912: data = 8'hf5;
      17'd70913: data = 8'h01;
      17'd70914: data = 8'hfc;
      17'd70915: data = 8'hf1;
      17'd70916: data = 8'h05;
      17'd70917: data = 8'h06;
      17'd70918: data = 8'hf4;
      17'd70919: data = 8'h0a;
      17'd70920: data = 8'h0d;
      17'd70921: data = 8'hfd;
      17'd70922: data = 8'h00;
      17'd70923: data = 8'h09;
      17'd70924: data = 8'hfd;
      17'd70925: data = 8'hef;
      17'd70926: data = 8'hfe;
      17'd70927: data = 8'hf9;
      17'd70928: data = 8'heb;
      17'd70929: data = 8'hfa;
      17'd70930: data = 8'hfc;
      17'd70931: data = 8'hf5;
      17'd70932: data = 8'hf5;
      17'd70933: data = 8'h04;
      17'd70934: data = 8'hef;
      17'd70935: data = 8'hf4;
      17'd70936: data = 8'h02;
      17'd70937: data = 8'hf6;
      17'd70938: data = 8'hfc;
      17'd70939: data = 8'h01;
      17'd70940: data = 8'hfa;
      17'd70941: data = 8'hf6;
      17'd70942: data = 8'hfc;
      17'd70943: data = 8'h00;
      17'd70944: data = 8'hf5;
      17'd70945: data = 8'hfe;
      17'd70946: data = 8'hfe;
      17'd70947: data = 8'he9;
      17'd70948: data = 8'hf9;
      17'd70949: data = 8'hf4;
      17'd70950: data = 8'hf6;
      17'd70951: data = 8'hfd;
      17'd70952: data = 8'hf5;
      17'd70953: data = 8'hfd;
      17'd70954: data = 8'hf5;
      17'd70955: data = 8'hf6;
      17'd70956: data = 8'hfc;
      17'd70957: data = 8'hf4;
      17'd70958: data = 8'hfa;
      17'd70959: data = 8'hfc;
      17'd70960: data = 8'hf6;
      17'd70961: data = 8'hf6;
      17'd70962: data = 8'hfd;
      17'd70963: data = 8'hf9;
      17'd70964: data = 8'hf6;
      17'd70965: data = 8'hf6;
      17'd70966: data = 8'hf5;
      17'd70967: data = 8'hfa;
      17'd70968: data = 8'hfa;
      17'd70969: data = 8'hfc;
      17'd70970: data = 8'h02;
      17'd70971: data = 8'hf9;
      17'd70972: data = 8'hf4;
      17'd70973: data = 8'hf9;
      17'd70974: data = 8'hf2;
      17'd70975: data = 8'hf2;
      17'd70976: data = 8'hed;
      17'd70977: data = 8'hfa;
      17'd70978: data = 8'hf5;
      17'd70979: data = 8'hf2;
      17'd70980: data = 8'hfe;
      17'd70981: data = 8'hf4;
      17'd70982: data = 8'hf6;
      17'd70983: data = 8'hf4;
      17'd70984: data = 8'hf1;
      17'd70985: data = 8'hf5;
      17'd70986: data = 8'hf5;
      17'd70987: data = 8'hfa;
      17'd70988: data = 8'hf6;
      17'd70989: data = 8'hfa;
      17'd70990: data = 8'hfe;
      17'd70991: data = 8'hf2;
      17'd70992: data = 8'hf1;
      17'd70993: data = 8'hf5;
      17'd70994: data = 8'hf4;
      17'd70995: data = 8'hf9;
      17'd70996: data = 8'h00;
      17'd70997: data = 8'h02;
      17'd70998: data = 8'h00;
      17'd70999: data = 8'hfe;
      17'd71000: data = 8'hfe;
      17'd71001: data = 8'hfc;
      17'd71002: data = 8'hf9;
      17'd71003: data = 8'hfd;
      17'd71004: data = 8'hfd;
      17'd71005: data = 8'hfd;
      17'd71006: data = 8'h05;
      17'd71007: data = 8'h01;
      17'd71008: data = 8'hfc;
      17'd71009: data = 8'h04;
      17'd71010: data = 8'h00;
      17'd71011: data = 8'hfa;
      17'd71012: data = 8'hfe;
      17'd71013: data = 8'h01;
      17'd71014: data = 8'h05;
      17'd71015: data = 8'h00;
      17'd71016: data = 8'h04;
      17'd71017: data = 8'h05;
      17'd71018: data = 8'hfe;
      17'd71019: data = 8'hfe;
      17'd71020: data = 8'hfc;
      17'd71021: data = 8'h00;
      17'd71022: data = 8'h02;
      17'd71023: data = 8'h02;
      17'd71024: data = 8'h09;
      17'd71025: data = 8'h09;
      17'd71026: data = 8'h02;
      17'd71027: data = 8'h01;
      17'd71028: data = 8'h02;
      17'd71029: data = 8'h00;
      17'd71030: data = 8'hfe;
      17'd71031: data = 8'hfe;
      17'd71032: data = 8'hfc;
      17'd71033: data = 8'hfd;
      17'd71034: data = 8'h00;
      17'd71035: data = 8'hfc;
      17'd71036: data = 8'hf6;
      17'd71037: data = 8'hfc;
      17'd71038: data = 8'hf9;
      17'd71039: data = 8'hf2;
      17'd71040: data = 8'hfd;
      17'd71041: data = 8'h01;
      17'd71042: data = 8'hfd;
      17'd71043: data = 8'h02;
      17'd71044: data = 8'h04;
      17'd71045: data = 8'hfd;
      17'd71046: data = 8'hf6;
      17'd71047: data = 8'hfd;
      17'd71048: data = 8'hfe;
      17'd71049: data = 8'hfc;
      17'd71050: data = 8'h02;
      17'd71051: data = 8'h01;
      17'd71052: data = 8'hfc;
      17'd71053: data = 8'h00;
      17'd71054: data = 8'h00;
      17'd71055: data = 8'hfe;
      17'd71056: data = 8'h00;
      17'd71057: data = 8'h00;
      17'd71058: data = 8'h01;
      17'd71059: data = 8'h00;
      17'd71060: data = 8'h02;
      17'd71061: data = 8'h06;
      17'd71062: data = 8'h01;
      17'd71063: data = 8'h02;
      17'd71064: data = 8'h04;
      17'd71065: data = 8'h02;
      17'd71066: data = 8'h02;
      17'd71067: data = 8'h06;
      17'd71068: data = 8'h0a;
      17'd71069: data = 8'h02;
      17'd71070: data = 8'h04;
      17'd71071: data = 8'h0c;
      17'd71072: data = 8'h06;
      17'd71073: data = 8'h02;
      17'd71074: data = 8'h09;
      17'd71075: data = 8'h06;
      17'd71076: data = 8'h05;
      17'd71077: data = 8'h0a;
      17'd71078: data = 8'h0c;
      17'd71079: data = 8'h09;
      17'd71080: data = 8'h0a;
      17'd71081: data = 8'h0c;
      17'd71082: data = 8'h06;
      17'd71083: data = 8'h02;
      17'd71084: data = 8'h04;
      17'd71085: data = 8'h02;
      17'd71086: data = 8'hfe;
      17'd71087: data = 8'h04;
      17'd71088: data = 8'h05;
      17'd71089: data = 8'hfe;
      17'd71090: data = 8'h02;
      17'd71091: data = 8'h04;
      17'd71092: data = 8'h02;
      17'd71093: data = 8'h02;
      17'd71094: data = 8'h06;
      17'd71095: data = 8'h06;
      17'd71096: data = 8'h06;
      17'd71097: data = 8'h06;
      17'd71098: data = 8'h05;
      17'd71099: data = 8'h02;
      17'd71100: data = 8'h02;
      17'd71101: data = 8'h01;
      17'd71102: data = 8'h00;
      17'd71103: data = 8'h01;
      17'd71104: data = 8'h01;
      17'd71105: data = 8'hfe;
      17'd71106: data = 8'h01;
      17'd71107: data = 8'h05;
      17'd71108: data = 8'h01;
      17'd71109: data = 8'h01;
      17'd71110: data = 8'h00;
      17'd71111: data = 8'h00;
      17'd71112: data = 8'h01;
      17'd71113: data = 8'h05;
      17'd71114: data = 8'h05;
      17'd71115: data = 8'h05;
      17'd71116: data = 8'h02;
      17'd71117: data = 8'h00;
      17'd71118: data = 8'h00;
      17'd71119: data = 8'h00;
      17'd71120: data = 8'hfe;
      17'd71121: data = 8'h01;
      17'd71122: data = 8'h02;
      17'd71123: data = 8'h01;
      17'd71124: data = 8'h04;
      17'd71125: data = 8'h04;
      17'd71126: data = 8'h04;
      17'd71127: data = 8'h0a;
      17'd71128: data = 8'h0d;
      17'd71129: data = 8'h02;
      17'd71130: data = 8'hfd;
      17'd71131: data = 8'h05;
      17'd71132: data = 8'h0c;
      17'd71133: data = 8'h04;
      17'd71134: data = 8'h00;
      17'd71135: data = 8'hfe;
      17'd71136: data = 8'h04;
      17'd71137: data = 8'h04;
      17'd71138: data = 8'h00;
      17'd71139: data = 8'h00;
      17'd71140: data = 8'h04;
      17'd71141: data = 8'h0a;
      17'd71142: data = 8'h01;
      17'd71143: data = 8'hfc;
      17'd71144: data = 8'hfd;
      17'd71145: data = 8'h02;
      17'd71146: data = 8'h04;
      17'd71147: data = 8'hfe;
      17'd71148: data = 8'hfc;
      17'd71149: data = 8'hfe;
      17'd71150: data = 8'hfe;
      17'd71151: data = 8'h00;
      17'd71152: data = 8'h00;
      17'd71153: data = 8'hfd;
      17'd71154: data = 8'hfd;
      17'd71155: data = 8'h00;
      17'd71156: data = 8'h04;
      17'd71157: data = 8'h02;
      17'd71158: data = 8'h01;
      17'd71159: data = 8'h01;
      17'd71160: data = 8'h01;
      17'd71161: data = 8'h06;
      17'd71162: data = 8'h02;
      17'd71163: data = 8'hf9;
      17'd71164: data = 8'hfc;
      17'd71165: data = 8'hfe;
      17'd71166: data = 8'h00;
      17'd71167: data = 8'h00;
      17'd71168: data = 8'hfc;
      17'd71169: data = 8'hfd;
      17'd71170: data = 8'h04;
      17'd71171: data = 8'h01;
      17'd71172: data = 8'hfa;
      17'd71173: data = 8'hfc;
      17'd71174: data = 8'h05;
      17'd71175: data = 8'h06;
      17'd71176: data = 8'h01;
      17'd71177: data = 8'h01;
      17'd71178: data = 8'h00;
      17'd71179: data = 8'h00;
      17'd71180: data = 8'h05;
      17'd71181: data = 8'h01;
      17'd71182: data = 8'hfe;
      17'd71183: data = 8'h04;
      17'd71184: data = 8'h04;
      17'd71185: data = 8'h02;
      17'd71186: data = 8'h02;
      17'd71187: data = 8'h06;
      17'd71188: data = 8'h06;
      17'd71189: data = 8'h02;
      17'd71190: data = 8'h05;
      17'd71191: data = 8'h04;
      17'd71192: data = 8'hfe;
      17'd71193: data = 8'h02;
      17'd71194: data = 8'h02;
      17'd71195: data = 8'h01;
      17'd71196: data = 8'h04;
      17'd71197: data = 8'h01;
      17'd71198: data = 8'h00;
      17'd71199: data = 8'h01;
      17'd71200: data = 8'h04;
      17'd71201: data = 8'h05;
      17'd71202: data = 8'h02;
      17'd71203: data = 8'h01;
      17'd71204: data = 8'h02;
      17'd71205: data = 8'h02;
      17'd71206: data = 8'h01;
      17'd71207: data = 8'hfe;
      17'd71208: data = 8'h01;
      17'd71209: data = 8'h02;
      17'd71210: data = 8'h00;
      17'd71211: data = 8'h01;
      17'd71212: data = 8'h04;
      17'd71213: data = 8'hfe;
      17'd71214: data = 8'h04;
      17'd71215: data = 8'h09;
      17'd71216: data = 8'hfe;
      17'd71217: data = 8'h00;
      17'd71218: data = 8'hfe;
      17'd71219: data = 8'hfc;
      17'd71220: data = 8'hfa;
      17'd71221: data = 8'hf9;
      17'd71222: data = 8'hf9;
      17'd71223: data = 8'hfa;
      17'd71224: data = 8'hf5;
      17'd71225: data = 8'hfc;
      17'd71226: data = 8'hfa;
      17'd71227: data = 8'hf5;
      17'd71228: data = 8'hfe;
      17'd71229: data = 8'hfc;
      17'd71230: data = 8'hfa;
      17'd71231: data = 8'h00;
      17'd71232: data = 8'hfd;
      17'd71233: data = 8'hfd;
      17'd71234: data = 8'h01;
      17'd71235: data = 8'h00;
      17'd71236: data = 8'h00;
      17'd71237: data = 8'hfd;
      17'd71238: data = 8'h00;
      17'd71239: data = 8'h01;
      17'd71240: data = 8'hfd;
      17'd71241: data = 8'h01;
      17'd71242: data = 8'h02;
      17'd71243: data = 8'hfd;
      17'd71244: data = 8'h00;
      17'd71245: data = 8'hfd;
      17'd71246: data = 8'hfc;
      17'd71247: data = 8'hfd;
      17'd71248: data = 8'hf9;
      17'd71249: data = 8'hfa;
      17'd71250: data = 8'hf9;
      17'd71251: data = 8'hf5;
      17'd71252: data = 8'hfe;
      17'd71253: data = 8'hfc;
      17'd71254: data = 8'hf9;
      17'd71255: data = 8'hf9;
      17'd71256: data = 8'hf9;
      17'd71257: data = 8'hfd;
      17'd71258: data = 8'hfd;
      17'd71259: data = 8'hfc;
      17'd71260: data = 8'h00;
      17'd71261: data = 8'hfc;
      17'd71262: data = 8'hfc;
      17'd71263: data = 8'hfc;
      17'd71264: data = 8'hf2;
      17'd71265: data = 8'hf9;
      17'd71266: data = 8'hfc;
      17'd71267: data = 8'hf6;
      17'd71268: data = 8'hfa;
      17'd71269: data = 8'hfa;
      17'd71270: data = 8'hfa;
      17'd71271: data = 8'hfc;
      17'd71272: data = 8'hfa;
      17'd71273: data = 8'hfc;
      17'd71274: data = 8'hf6;
      17'd71275: data = 8'hf4;
      17'd71276: data = 8'hf6;
      17'd71277: data = 8'hfa;
      17'd71278: data = 8'hfc;
      17'd71279: data = 8'hfc;
      17'd71280: data = 8'hf9;
      17'd71281: data = 8'hfa;
      17'd71282: data = 8'hfc;
      17'd71283: data = 8'hf6;
      17'd71284: data = 8'hfd;
      17'd71285: data = 8'hfe;
      17'd71286: data = 8'h04;
      17'd71287: data = 8'h01;
      17'd71288: data = 8'hfa;
      17'd71289: data = 8'hfa;
      17'd71290: data = 8'hfc;
      17'd71291: data = 8'hf6;
      17'd71292: data = 8'hf9;
      17'd71293: data = 8'hf6;
      17'd71294: data = 8'hf9;
      17'd71295: data = 8'hfa;
      17'd71296: data = 8'hf9;
      17'd71297: data = 8'hfa;
      17'd71298: data = 8'hfd;
      17'd71299: data = 8'hfd;
      17'd71300: data = 8'hfc;
      17'd71301: data = 8'hfd;
      17'd71302: data = 8'h01;
      17'd71303: data = 8'hfe;
      17'd71304: data = 8'hfc;
      17'd71305: data = 8'hfe;
      17'd71306: data = 8'hfe;
      17'd71307: data = 8'hf9;
      17'd71308: data = 8'hf4;
      17'd71309: data = 8'hf5;
      17'd71310: data = 8'hf4;
      17'd71311: data = 8'hf5;
      17'd71312: data = 8'hf9;
      17'd71313: data = 8'hfa;
      17'd71314: data = 8'hfd;
      17'd71315: data = 8'h00;
      17'd71316: data = 8'hfe;
      17'd71317: data = 8'hfd;
      17'd71318: data = 8'hfe;
      17'd71319: data = 8'h01;
      17'd71320: data = 8'hfc;
      17'd71321: data = 8'hf9;
      17'd71322: data = 8'hfe;
      17'd71323: data = 8'hfc;
      17'd71324: data = 8'hf9;
      17'd71325: data = 8'hfc;
      17'd71326: data = 8'hfe;
      17'd71327: data = 8'hfa;
      17'd71328: data = 8'hfa;
      17'd71329: data = 8'h04;
      17'd71330: data = 8'h01;
      17'd71331: data = 8'h01;
      17'd71332: data = 8'h05;
      17'd71333: data = 8'h00;
      17'd71334: data = 8'h01;
      17'd71335: data = 8'h04;
      17'd71336: data = 8'hfe;
      17'd71337: data = 8'hf9;
      17'd71338: data = 8'hfa;
      17'd71339: data = 8'hfc;
      17'd71340: data = 8'hf6;
      17'd71341: data = 8'hf9;
      17'd71342: data = 8'hfe;
      17'd71343: data = 8'hfd;
      17'd71344: data = 8'hfa;
      17'd71345: data = 8'h02;
      17'd71346: data = 8'h00;
      17'd71347: data = 8'hfc;
      17'd71348: data = 8'h01;
      17'd71349: data = 8'h00;
      17'd71350: data = 8'h00;
      17'd71351: data = 8'h02;
      17'd71352: data = 8'hfe;
      17'd71353: data = 8'h00;
      17'd71354: data = 8'h02;
      17'd71355: data = 8'h00;
      17'd71356: data = 8'h00;
      17'd71357: data = 8'h01;
      17'd71358: data = 8'h01;
      17'd71359: data = 8'h01;
      17'd71360: data = 8'h02;
      17'd71361: data = 8'h05;
      17'd71362: data = 8'h02;
      17'd71363: data = 8'h00;
      17'd71364: data = 8'h04;
      17'd71365: data = 8'h00;
      17'd71366: data = 8'h01;
      17'd71367: data = 8'h04;
      17'd71368: data = 8'hfe;
      17'd71369: data = 8'h00;
      17'd71370: data = 8'h04;
      17'd71371: data = 8'hfe;
      17'd71372: data = 8'h00;
      17'd71373: data = 8'h05;
      17'd71374: data = 8'h04;
      17'd71375: data = 8'h02;
      17'd71376: data = 8'h04;
      17'd71377: data = 8'h09;
      17'd71378: data = 8'h06;
      17'd71379: data = 8'h09;
      17'd71380: data = 8'h0d;
      17'd71381: data = 8'h05;
      17'd71382: data = 8'h06;
      17'd71383: data = 8'h0a;
      17'd71384: data = 8'h04;
      17'd71385: data = 8'h04;
      17'd71386: data = 8'h05;
      17'd71387: data = 8'h04;
      17'd71388: data = 8'h05;
      17'd71389: data = 8'h06;
      17'd71390: data = 8'h05;
      17'd71391: data = 8'h02;
      17'd71392: data = 8'h04;
      17'd71393: data = 8'h09;
      17'd71394: data = 8'h05;
      17'd71395: data = 8'h01;
      17'd71396: data = 8'h01;
      17'd71397: data = 8'h00;
      17'd71398: data = 8'h00;
      17'd71399: data = 8'h01;
      17'd71400: data = 8'h00;
      17'd71401: data = 8'hfe;
      17'd71402: data = 8'hfe;
      17'd71403: data = 8'h01;
      17'd71404: data = 8'h02;
      17'd71405: data = 8'h02;
      17'd71406: data = 8'h04;
      17'd71407: data = 8'h05;
      17'd71408: data = 8'h05;
      17'd71409: data = 8'h04;
      17'd71410: data = 8'h02;
      17'd71411: data = 8'h00;
      17'd71412: data = 8'h00;
      17'd71413: data = 8'h00;
      17'd71414: data = 8'h00;
      17'd71415: data = 8'hfd;
      17'd71416: data = 8'hf9;
      17'd71417: data = 8'hf6;
      17'd71418: data = 8'hfa;
      17'd71419: data = 8'hfe;
      17'd71420: data = 8'h00;
      17'd71421: data = 8'h02;
      17'd71422: data = 8'h02;
      17'd71423: data = 8'h05;
      17'd71424: data = 8'h0a;
      17'd71425: data = 8'h0a;
      17'd71426: data = 8'h09;
      17'd71427: data = 8'h06;
      17'd71428: data = 8'h06;
      17'd71429: data = 8'h06;
      17'd71430: data = 8'h04;
      17'd71431: data = 8'hfe;
      17'd71432: data = 8'hfe;
      17'd71433: data = 8'hfe;
      17'd71434: data = 8'h00;
      17'd71435: data = 8'h00;
      17'd71436: data = 8'hfe;
      17'd71437: data = 8'h00;
      17'd71438: data = 8'h01;
      17'd71439: data = 8'h02;
      17'd71440: data = 8'h05;
      17'd71441: data = 8'h06;
      17'd71442: data = 8'h05;
      17'd71443: data = 8'h05;
      17'd71444: data = 8'h06;
      17'd71445: data = 8'h05;
      17'd71446: data = 8'h02;
      17'd71447: data = 8'h01;
      17'd71448: data = 8'h01;
      17'd71449: data = 8'h00;
      17'd71450: data = 8'h00;
      17'd71451: data = 8'h00;
      17'd71452: data = 8'hfd;
      17'd71453: data = 8'hfd;
      17'd71454: data = 8'h00;
      17'd71455: data = 8'h00;
      17'd71456: data = 8'h00;
      17'd71457: data = 8'h01;
      17'd71458: data = 8'hfe;
      17'd71459: data = 8'hfe;
      17'd71460: data = 8'h00;
      17'd71461: data = 8'hfd;
      17'd71462: data = 8'hf9;
      17'd71463: data = 8'hf9;
      17'd71464: data = 8'hfa;
      17'd71465: data = 8'hfa;
      17'd71466: data = 8'hfa;
      17'd71467: data = 8'hfa;
      17'd71468: data = 8'hfd;
      17'd71469: data = 8'hfc;
      17'd71470: data = 8'hfd;
      17'd71471: data = 8'h00;
      17'd71472: data = 8'h00;
      17'd71473: data = 8'h02;
      17'd71474: data = 8'h04;
      17'd71475: data = 8'h04;
      17'd71476: data = 8'h0a;
      17'd71477: data = 8'h09;
      17'd71478: data = 8'h05;
      17'd71479: data = 8'h06;
      17'd71480: data = 8'h05;
      17'd71481: data = 8'h02;
      17'd71482: data = 8'h02;
      17'd71483: data = 8'h01;
      17'd71484: data = 8'h01;
      17'd71485: data = 8'h04;
      17'd71486: data = 8'h02;
      17'd71487: data = 8'h04;
      17'd71488: data = 8'h01;
      17'd71489: data = 8'h01;
      17'd71490: data = 8'h01;
      17'd71491: data = 8'h00;
      17'd71492: data = 8'h01;
      17'd71493: data = 8'h00;
      17'd71494: data = 8'hfe;
      17'd71495: data = 8'hfc;
      17'd71496: data = 8'hfc;
      17'd71497: data = 8'hfc;
      17'd71498: data = 8'hfe;
      17'd71499: data = 8'hfd;
      17'd71500: data = 8'hfa;
      17'd71501: data = 8'hfe;
      17'd71502: data = 8'hfd;
      17'd71503: data = 8'h00;
      17'd71504: data = 8'h00;
      17'd71505: data = 8'hfe;
      17'd71506: data = 8'hfe;
      17'd71507: data = 8'hfd;
      17'd71508: data = 8'hfc;
      17'd71509: data = 8'hfa;
      17'd71510: data = 8'hf6;
      17'd71511: data = 8'hf5;
      17'd71512: data = 8'hf6;
      17'd71513: data = 8'hf9;
      17'd71514: data = 8'hf6;
      17'd71515: data = 8'hf5;
      17'd71516: data = 8'hf6;
      17'd71517: data = 8'hfa;
      17'd71518: data = 8'hfc;
      17'd71519: data = 8'hfc;
      17'd71520: data = 8'hfe;
      17'd71521: data = 8'hfd;
      17'd71522: data = 8'hfe;
      17'd71523: data = 8'h01;
      17'd71524: data = 8'h00;
      17'd71525: data = 8'hfd;
      17'd71526: data = 8'hfc;
      17'd71527: data = 8'hfd;
      17'd71528: data = 8'hfd;
      17'd71529: data = 8'hfd;
      17'd71530: data = 8'hfe;
      17'd71531: data = 8'hfc;
      17'd71532: data = 8'hfe;
      17'd71533: data = 8'h01;
      17'd71534: data = 8'hfe;
      17'd71535: data = 8'hfe;
      17'd71536: data = 8'hfd;
      17'd71537: data = 8'hfd;
      17'd71538: data = 8'hfe;
      17'd71539: data = 8'h00;
      17'd71540: data = 8'hfd;
      17'd71541: data = 8'hfa;
      17'd71542: data = 8'hfc;
      17'd71543: data = 8'hfc;
      17'd71544: data = 8'hfd;
      17'd71545: data = 8'hfa;
      17'd71546: data = 8'hfc;
      17'd71547: data = 8'hfd;
      17'd71548: data = 8'hfd;
      17'd71549: data = 8'h01;
      17'd71550: data = 8'h01;
      17'd71551: data = 8'h02;
      17'd71552: data = 8'h02;
      17'd71553: data = 8'h02;
      17'd71554: data = 8'h02;
      17'd71555: data = 8'h00;
      17'd71556: data = 8'hfe;
      17'd71557: data = 8'hfd;
      17'd71558: data = 8'hfe;
      17'd71559: data = 8'hfe;
      17'd71560: data = 8'hfd;
      17'd71561: data = 8'hfd;
      17'd71562: data = 8'hfa;
      17'd71563: data = 8'hfc;
      17'd71564: data = 8'hfe;
      17'd71565: data = 8'hfc;
      17'd71566: data = 8'hfd;
      17'd71567: data = 8'hfd;
      17'd71568: data = 8'hfd;
      17'd71569: data = 8'hfd;
      17'd71570: data = 8'hfa;
      17'd71571: data = 8'hfa;
      17'd71572: data = 8'hf6;
      17'd71573: data = 8'hf9;
      17'd71574: data = 8'hf9;
      17'd71575: data = 8'hf5;
      17'd71576: data = 8'hfa;
      17'd71577: data = 8'hfd;
      17'd71578: data = 8'hfc;
      17'd71579: data = 8'hfc;
      17'd71580: data = 8'hfd;
      17'd71581: data = 8'hfd;
      17'd71582: data = 8'hfe;
      17'd71583: data = 8'hfd;
      17'd71584: data = 8'hfc;
      17'd71585: data = 8'hfc;
      17'd71586: data = 8'hfc;
      17'd71587: data = 8'hfc;
      17'd71588: data = 8'hfc;
      17'd71589: data = 8'hfc;
      17'd71590: data = 8'hfe;
      17'd71591: data = 8'hfe;
      17'd71592: data = 8'hfe;
      17'd71593: data = 8'hfd;
      17'd71594: data = 8'hfd;
      17'd71595: data = 8'h00;
      17'd71596: data = 8'hfe;
      17'd71597: data = 8'hfe;
      17'd71598: data = 8'hfd;
      17'd71599: data = 8'hfa;
      17'd71600: data = 8'hfc;
      17'd71601: data = 8'hfe;
      17'd71602: data = 8'hfd;
      17'd71603: data = 8'hfd;
      17'd71604: data = 8'hfe;
      17'd71605: data = 8'hfe;
      17'd71606: data = 8'h01;
      17'd71607: data = 8'h02;
      17'd71608: data = 8'h01;
      17'd71609: data = 8'h00;
      17'd71610: data = 8'h01;
      17'd71611: data = 8'h01;
      17'd71612: data = 8'h00;
      17'd71613: data = 8'h00;
      17'd71614: data = 8'hfd;
      17'd71615: data = 8'hfc;
      17'd71616: data = 8'hfc;
      17'd71617: data = 8'hfd;
      17'd71618: data = 8'hfc;
      17'd71619: data = 8'hfd;
      17'd71620: data = 8'hfe;
      17'd71621: data = 8'hfe;
      17'd71622: data = 8'h00;
      17'd71623: data = 8'h01;
      17'd71624: data = 8'h00;
      17'd71625: data = 8'h01;
      17'd71626: data = 8'h04;
      17'd71627: data = 8'h05;
      17'd71628: data = 8'h04;
      17'd71629: data = 8'h04;
      17'd71630: data = 8'h04;
      17'd71631: data = 8'h02;
      17'd71632: data = 8'h02;
      17'd71633: data = 8'h01;
      17'd71634: data = 8'h01;
      17'd71635: data = 8'h02;
      17'd71636: data = 8'h02;
      17'd71637: data = 8'h04;
      17'd71638: data = 8'h04;
      17'd71639: data = 8'h05;
      17'd71640: data = 8'h05;
      17'd71641: data = 8'h05;
      17'd71642: data = 8'h04;
      17'd71643: data = 8'h06;
      17'd71644: data = 8'h05;
      17'd71645: data = 8'h01;
      17'd71646: data = 8'h01;
      17'd71647: data = 8'h00;
      17'd71648: data = 8'h00;
      17'd71649: data = 8'h00;
      17'd71650: data = 8'h00;
      17'd71651: data = 8'hfe;
      17'd71652: data = 8'hfe;
      17'd71653: data = 8'h01;
      17'd71654: data = 8'h00;
      17'd71655: data = 8'h00;
      17'd71656: data = 8'h01;
      17'd71657: data = 8'h01;
      17'd71658: data = 8'h01;
      17'd71659: data = 8'hfe;
      17'd71660: data = 8'h00;
      17'd71661: data = 8'h01;
      17'd71662: data = 8'hfe;
      17'd71663: data = 8'hfe;
      17'd71664: data = 8'hfe;
      17'd71665: data = 8'h00;
      17'd71666: data = 8'hfe;
      17'd71667: data = 8'h00;
      17'd71668: data = 8'h01;
      17'd71669: data = 8'h02;
      17'd71670: data = 8'h04;
      17'd71671: data = 8'h02;
      17'd71672: data = 8'h02;
      17'd71673: data = 8'h02;
      17'd71674: data = 8'h02;
      17'd71675: data = 8'h01;
      17'd71676: data = 8'h01;
      17'd71677: data = 8'h01;
      17'd71678: data = 8'h00;
      17'd71679: data = 8'h01;
      17'd71680: data = 8'h02;
      17'd71681: data = 8'h02;
      17'd71682: data = 8'h01;
      17'd71683: data = 8'h02;
      17'd71684: data = 8'h04;
      17'd71685: data = 8'h05;
      17'd71686: data = 8'h06;
      17'd71687: data = 8'h05;
      17'd71688: data = 8'h04;
      17'd71689: data = 8'h05;
      17'd71690: data = 8'h05;
      17'd71691: data = 8'h01;
      17'd71692: data = 8'h02;
      17'd71693: data = 8'h02;
      17'd71694: data = 8'h01;
      17'd71695: data = 8'h02;
      17'd71696: data = 8'h00;
      17'd71697: data = 8'h00;
      17'd71698: data = 8'h00;
      17'd71699: data = 8'h00;
      17'd71700: data = 8'h00;
      17'd71701: data = 8'h00;
      17'd71702: data = 8'hfe;
      17'd71703: data = 8'hfe;
      17'd71704: data = 8'hfd;
      17'd71705: data = 8'hfe;
      17'd71706: data = 8'hfe;
      17'd71707: data = 8'hfe;
      17'd71708: data = 8'hfe;
      17'd71709: data = 8'hfa;
      17'd71710: data = 8'hfa;
      17'd71711: data = 8'hfc;
      17'd71712: data = 8'hfc;
      17'd71713: data = 8'hfc;
      17'd71714: data = 8'hfd;
      17'd71715: data = 8'hfe;
      17'd71716: data = 8'hfe;
      17'd71717: data = 8'hfe;
      17'd71718: data = 8'hfe;
      17'd71719: data = 8'hfd;
      17'd71720: data = 8'h00;
      17'd71721: data = 8'h01;
      17'd71722: data = 8'h02;
      17'd71723: data = 8'h00;
      17'd71724: data = 8'h00;
      17'd71725: data = 8'h00;
      17'd71726: data = 8'hfe;
      17'd71727: data = 8'hfe;
      17'd71728: data = 8'hfd;
      17'd71729: data = 8'hfd;
      17'd71730: data = 8'hfe;
      17'd71731: data = 8'h01;
      17'd71732: data = 8'h02;
      17'd71733: data = 8'h02;
      17'd71734: data = 8'h02;
      17'd71735: data = 8'h02;
      17'd71736: data = 8'h02;
      17'd71737: data = 8'h00;
      17'd71738: data = 8'h01;
      17'd71739: data = 8'h00;
      17'd71740: data = 8'h00;
      17'd71741: data = 8'h00;
      17'd71742: data = 8'h01;
      17'd71743: data = 8'h01;
      17'd71744: data = 8'h02;
      17'd71745: data = 8'h02;
      17'd71746: data = 8'h01;
      17'd71747: data = 8'h02;
      17'd71748: data = 8'h02;
      17'd71749: data = 8'h01;
      17'd71750: data = 8'h02;
      17'd71751: data = 8'h04;
      17'd71752: data = 8'h01;
      17'd71753: data = 8'h01;
      17'd71754: data = 8'h01;
      17'd71755: data = 8'hfe;
      17'd71756: data = 8'hfd;
      17'd71757: data = 8'h00;
      17'd71758: data = 8'hfe;
      17'd71759: data = 8'hfe;
      17'd71760: data = 8'hfe;
      17'd71761: data = 8'hfe;
      17'd71762: data = 8'hfd;
      17'd71763: data = 8'hfc;
      17'd71764: data = 8'hfc;
      17'd71765: data = 8'hfd;
      17'd71766: data = 8'hfe;
      17'd71767: data = 8'hfd;
      17'd71768: data = 8'hfe;
      17'd71769: data = 8'hfd;
      17'd71770: data = 8'hfc;
      17'd71771: data = 8'hfe;
      17'd71772: data = 8'hfe;
      17'd71773: data = 8'hfd;
      17'd71774: data = 8'hfd;
      17'd71775: data = 8'hfc;
      17'd71776: data = 8'hfc;
      17'd71777: data = 8'hfc;
      17'd71778: data = 8'hfd;
      17'd71779: data = 8'hfd;
      17'd71780: data = 8'h01;
      17'd71781: data = 8'h01;
      17'd71782: data = 8'h01;
      17'd71783: data = 8'h02;
      17'd71784: data = 8'h01;
      17'd71785: data = 8'h01;
      17'd71786: data = 8'h00;
      17'd71787: data = 8'h00;
      17'd71788: data = 8'h00;
      17'd71789: data = 8'hfd;
      17'd71790: data = 8'hfe;
      17'd71791: data = 8'hfe;
      17'd71792: data = 8'hfe;
      17'd71793: data = 8'hfe;
      17'd71794: data = 8'h00;
      17'd71795: data = 8'h00;
      17'd71796: data = 8'h00;
      17'd71797: data = 8'h00;
      17'd71798: data = 8'h01;
      17'd71799: data = 8'h00;
      17'd71800: data = 8'hfe;
      17'd71801: data = 8'hfe;
      17'd71802: data = 8'hfc;
      17'd71803: data = 8'hf9;
      17'd71804: data = 8'hfa;
      17'd71805: data = 8'hfc;
      17'd71806: data = 8'hf9;
      17'd71807: data = 8'hf6;
      17'd71808: data = 8'hfa;
      17'd71809: data = 8'hfa;
      17'd71810: data = 8'hfa;
      17'd71811: data = 8'hfa;
      17'd71812: data = 8'hf9;
      17'd71813: data = 8'hf9;
      17'd71814: data = 8'hf9;
      17'd71815: data = 8'hf9;
      17'd71816: data = 8'hf9;
      17'd71817: data = 8'hfc;
      17'd71818: data = 8'hfc;
      17'd71819: data = 8'hfa;
      17'd71820: data = 8'hfc;
      17'd71821: data = 8'hfc;
      17'd71822: data = 8'hf9;
      17'd71823: data = 8'hfa;
      17'd71824: data = 8'hfc;
      17'd71825: data = 8'hfc;
      17'd71826: data = 8'hfd;
      17'd71827: data = 8'hfd;
      17'd71828: data = 8'hfd;
      17'd71829: data = 8'hfd;
      17'd71830: data = 8'hfe;
      17'd71831: data = 8'hfe;
      17'd71832: data = 8'hfe;
      17'd71833: data = 8'h00;
      17'd71834: data = 8'h01;
      17'd71835: data = 8'h01;
      17'd71836: data = 8'h02;
      17'd71837: data = 8'h01;
      17'd71838: data = 8'hfe;
      17'd71839: data = 8'h00;
      17'd71840: data = 8'h00;
      17'd71841: data = 8'hfe;
      17'd71842: data = 8'hfe;
      17'd71843: data = 8'hfe;
      17'd71844: data = 8'hfe;
      17'd71845: data = 8'hfe;
      17'd71846: data = 8'hfe;
      17'd71847: data = 8'hfe;
      17'd71848: data = 8'h00;
      17'd71849: data = 8'h00;
      17'd71850: data = 8'hfe;
      17'd71851: data = 8'hfc;
      17'd71852: data = 8'hfc;
      17'd71853: data = 8'hfd;
      17'd71854: data = 8'hfc;
      17'd71855: data = 8'hfd;
      17'd71856: data = 8'hfd;
      17'd71857: data = 8'hfd;
      17'd71858: data = 8'hfd;
      17'd71859: data = 8'hf9;
      17'd71860: data = 8'hfc;
      17'd71861: data = 8'hfd;
      17'd71862: data = 8'hfd;
      17'd71863: data = 8'hfd;
      17'd71864: data = 8'hfe;
      17'd71865: data = 8'hfe;
      17'd71866: data = 8'hfe;
      17'd71867: data = 8'hfe;
      17'd71868: data = 8'hfe;
      17'd71869: data = 8'h00;
      17'd71870: data = 8'h01;
      17'd71871: data = 8'h01;
      17'd71872: data = 8'h00;
      17'd71873: data = 8'h00;
      17'd71874: data = 8'h01;
      17'd71875: data = 8'h00;
      17'd71876: data = 8'h01;
      17'd71877: data = 8'h01;
      17'd71878: data = 8'hfd;
      17'd71879: data = 8'hfe;
      17'd71880: data = 8'hfd;
      17'd71881: data = 8'hfe;
      17'd71882: data = 8'h00;
      17'd71883: data = 8'hfe;
      17'd71884: data = 8'h01;
      17'd71885: data = 8'h00;
      17'd71886: data = 8'h00;
      17'd71887: data = 8'hfe;
      17'd71888: data = 8'hfc;
      17'd71889: data = 8'hfa;
      17'd71890: data = 8'hfa;
      17'd71891: data = 8'hfc;
      17'd71892: data = 8'hf9;
      17'd71893: data = 8'hf9;
      17'd71894: data = 8'hf9;
      17'd71895: data = 8'hfa;
      17'd71896: data = 8'hfc;
      17'd71897: data = 8'hfa;
      17'd71898: data = 8'hfc;
      17'd71899: data = 8'hfc;
      17'd71900: data = 8'hfd;
      17'd71901: data = 8'hfe;
      17'd71902: data = 8'hfc;
      17'd71903: data = 8'hfd;
      17'd71904: data = 8'hfd;
      17'd71905: data = 8'hfd;
      17'd71906: data = 8'hfd;
      17'd71907: data = 8'hfd;
      17'd71908: data = 8'h00;
      17'd71909: data = 8'h01;
      17'd71910: data = 8'h00;
      17'd71911: data = 8'h02;
      17'd71912: data = 8'h02;
      17'd71913: data = 8'h00;
      17'd71914: data = 8'h01;
      17'd71915: data = 8'h01;
      17'd71916: data = 8'h01;
      17'd71917: data = 8'h01;
      17'd71918: data = 8'h02;
      17'd71919: data = 8'h04;
      17'd71920: data = 8'h04;
      17'd71921: data = 8'h04;
      17'd71922: data = 8'h04;
      17'd71923: data = 8'h05;
      17'd71924: data = 8'h02;
      17'd71925: data = 8'h01;
      17'd71926: data = 8'h01;
      17'd71927: data = 8'h01;
      17'd71928: data = 8'h01;
      17'd71929: data = 8'h02;
      17'd71930: data = 8'h01;
      17'd71931: data = 8'h02;
      17'd71932: data = 8'h01;
      17'd71933: data = 8'hfe;
      17'd71934: data = 8'h00;
      17'd71935: data = 8'h01;
      17'd71936: data = 8'h01;
      17'd71937: data = 8'h01;
      17'd71938: data = 8'h00;
      17'd71939: data = 8'h01;
      17'd71940: data = 8'h01;
      17'd71941: data = 8'hfd;
      17'd71942: data = 8'hfc;
      17'd71943: data = 8'hfd;
      17'd71944: data = 8'hfd;
      17'd71945: data = 8'hfe;
      17'd71946: data = 8'hfd;
      17'd71947: data = 8'hfe;
      17'd71948: data = 8'h00;
      17'd71949: data = 8'hfe;
      17'd71950: data = 8'hfd;
      17'd71951: data = 8'hfe;
      17'd71952: data = 8'hfe;
      17'd71953: data = 8'h00;
      17'd71954: data = 8'hfd;
      17'd71955: data = 8'hfe;
      17'd71956: data = 8'h00;
      17'd71957: data = 8'h00;
      17'd71958: data = 8'h00;
      17'd71959: data = 8'h00;
      17'd71960: data = 8'h00;
      17'd71961: data = 8'h01;
      17'd71962: data = 8'h00;
      17'd71963: data = 8'h01;
      17'd71964: data = 8'h02;
      17'd71965: data = 8'h01;
      17'd71966: data = 8'h02;
      17'd71967: data = 8'h04;
      17'd71968: data = 8'h04;
      17'd71969: data = 8'h04;
      17'd71970: data = 8'h02;
      17'd71971: data = 8'h04;
      17'd71972: data = 8'h05;
      17'd71973: data = 8'h04;
      17'd71974: data = 8'h04;
      17'd71975: data = 8'h02;
      17'd71976: data = 8'h04;
      17'd71977: data = 8'h05;
      17'd71978: data = 8'h02;
      17'd71979: data = 8'h02;
      17'd71980: data = 8'h02;
      17'd71981: data = 8'h05;
      17'd71982: data = 8'h04;
      17'd71983: data = 8'h02;
      17'd71984: data = 8'h04;
      17'd71985: data = 8'h02;
      17'd71986: data = 8'h02;
      17'd71987: data = 8'h01;
      17'd71988: data = 8'h01;
      17'd71989: data = 8'h01;
      17'd71990: data = 8'hfe;
      17'd71991: data = 8'h00;
      17'd71992: data = 8'h00;
      17'd71993: data = 8'hfc;
      17'd71994: data = 8'hfe;
      17'd71995: data = 8'h00;
      17'd71996: data = 8'hfe;
      17'd71997: data = 8'hfe;
      17'd71998: data = 8'hfe;
      17'd71999: data = 8'hfe;
      17'd72000: data = 8'h00;
      17'd72001: data = 8'hfe;
      17'd72002: data = 8'hfd;
      17'd72003: data = 8'hfd;
      17'd72004: data = 8'hfd;
      17'd72005: data = 8'hfd;
      17'd72006: data = 8'hfd;
      17'd72007: data = 8'hfe;
      17'd72008: data = 8'hfe;
      17'd72009: data = 8'hfd;
      17'd72010: data = 8'hfd;
      17'd72011: data = 8'h00;
      17'd72012: data = 8'h00;
      17'd72013: data = 8'h00;
      17'd72014: data = 8'h00;
      17'd72015: data = 8'h00;
      17'd72016: data = 8'h00;
      17'd72017: data = 8'h01;
      17'd72018: data = 8'h01;
      17'd72019: data = 8'h02;
      17'd72020: data = 8'h01;
      17'd72021: data = 8'h01;
      17'd72022: data = 8'h02;
      17'd72023: data = 8'h01;
      17'd72024: data = 8'h02;
      17'd72025: data = 8'h04;
      17'd72026: data = 8'h02;
      17'd72027: data = 8'h02;
      17'd72028: data = 8'h02;
      17'd72029: data = 8'h04;
      17'd72030: data = 8'h02;
      17'd72031: data = 8'h01;
      17'd72032: data = 8'h02;
      17'd72033: data = 8'h04;
      17'd72034: data = 8'h01;
      17'd72035: data = 8'h00;
      17'd72036: data = 8'h00;
      17'd72037: data = 8'h00;
      17'd72038: data = 8'hfe;
      17'd72039: data = 8'hfe;
      17'd72040: data = 8'hfd;
      17'd72041: data = 8'hfc;
      17'd72042: data = 8'hfd;
      17'd72043: data = 8'hfd;
      17'd72044: data = 8'hfc;
      17'd72045: data = 8'hfa;
      17'd72046: data = 8'hfc;
      17'd72047: data = 8'hfc;
      17'd72048: data = 8'hfd;
      17'd72049: data = 8'hfd;
      17'd72050: data = 8'hfc;
      17'd72051: data = 8'hfd;
      17'd72052: data = 8'hfe;
      17'd72053: data = 8'hfe;
      17'd72054: data = 8'hfd;
      17'd72055: data = 8'hfd;
      17'd72056: data = 8'hfc;
      17'd72057: data = 8'hfc;
      17'd72058: data = 8'hfa;
      17'd72059: data = 8'hfc;
      17'd72060: data = 8'hfc;
      17'd72061: data = 8'hfd;
      17'd72062: data = 8'hfe;
      17'd72063: data = 8'hfe;
      17'd72064: data = 8'h00;
      17'd72065: data = 8'hfe;
      17'd72066: data = 8'h00;
      17'd72067: data = 8'h00;
      17'd72068: data = 8'h00;
      17'd72069: data = 8'hfd;
      17'd72070: data = 8'hfe;
      17'd72071: data = 8'h00;
      17'd72072: data = 8'hfe;
      17'd72073: data = 8'hfd;
      17'd72074: data = 8'hfe;
      17'd72075: data = 8'hfe;
      17'd72076: data = 8'hfe;
      17'd72077: data = 8'hfe;
      17'd72078: data = 8'hfd;
      17'd72079: data = 8'hfd;
      17'd72080: data = 8'hfd;
      17'd72081: data = 8'hfd;
      17'd72082: data = 8'hfd;
      17'd72083: data = 8'hfe;
      17'd72084: data = 8'hfd;
      17'd72085: data = 8'hfe;
      17'd72086: data = 8'hfd;
      17'd72087: data = 8'hfd;
      17'd72088: data = 8'hfd;
      17'd72089: data = 8'hfc;
      17'd72090: data = 8'hfc;
      17'd72091: data = 8'hfc;
      17'd72092: data = 8'hfd;
      17'd72093: data = 8'hfd;
      17'd72094: data = 8'hfc;
      17'd72095: data = 8'hfd;
      17'd72096: data = 8'hfd;
      17'd72097: data = 8'hfd;
      17'd72098: data = 8'h00;
      17'd72099: data = 8'hfe;
      17'd72100: data = 8'hfe;
      17'd72101: data = 8'h00;
      17'd72102: data = 8'hfe;
      17'd72103: data = 8'h00;
      17'd72104: data = 8'h02;
      17'd72105: data = 8'h02;
      17'd72106: data = 8'h02;
      17'd72107: data = 8'h01;
      17'd72108: data = 8'hfe;
      17'd72109: data = 8'h01;
      17'd72110: data = 8'h02;
      17'd72111: data = 8'h01;
      17'd72112: data = 8'h02;
      17'd72113: data = 8'h01;
      17'd72114: data = 8'h02;
      17'd72115: data = 8'h01;
      17'd72116: data = 8'h00;
      17'd72117: data = 8'h01;
      17'd72118: data = 8'h00;
      17'd72119: data = 8'h01;
      17'd72120: data = 8'h01;
      17'd72121: data = 8'h00;
      17'd72122: data = 8'h00;
      17'd72123: data = 8'hfe;
      17'd72124: data = 8'hfe;
      17'd72125: data = 8'h00;
      17'd72126: data = 8'hfd;
      17'd72127: data = 8'hfe;
      17'd72128: data = 8'hfe;
      17'd72129: data = 8'hfe;
      17'd72130: data = 8'h00;
      17'd72131: data = 8'h00;
      17'd72132: data = 8'hfd;
      17'd72133: data = 8'hfd;
      17'd72134: data = 8'hfc;
      17'd72135: data = 8'hfe;
      17'd72136: data = 8'hfd;
      17'd72137: data = 8'hfd;
      17'd72138: data = 8'hfe;
      17'd72139: data = 8'hfc;
      17'd72140: data = 8'hfc;
      17'd72141: data = 8'hfd;
      17'd72142: data = 8'hfd;
      17'd72143: data = 8'hfe;
      17'd72144: data = 8'h01;
      17'd72145: data = 8'h00;
      17'd72146: data = 8'h00;
      17'd72147: data = 8'h01;
      17'd72148: data = 8'h00;
      17'd72149: data = 8'h00;
      17'd72150: data = 8'h00;
      17'd72151: data = 8'h00;
      17'd72152: data = 8'h00;
      17'd72153: data = 8'h01;
      17'd72154: data = 8'hfe;
      17'd72155: data = 8'hfe;
      17'd72156: data = 8'h00;
      17'd72157: data = 8'hfe;
      17'd72158: data = 8'h02;
      17'd72159: data = 8'h02;
      17'd72160: data = 8'h02;
      17'd72161: data = 8'h02;
      17'd72162: data = 8'h01;
      17'd72163: data = 8'h01;
      17'd72164: data = 8'h00;
      17'd72165: data = 8'h00;
      17'd72166: data = 8'hfd;
      17'd72167: data = 8'hfe;
      17'd72168: data = 8'hfd;
      17'd72169: data = 8'hfa;
      17'd72170: data = 8'hfc;
      17'd72171: data = 8'hfc;
      17'd72172: data = 8'hfa;
      17'd72173: data = 8'hfa;
      17'd72174: data = 8'hfd;
      17'd72175: data = 8'hfe;
      17'd72176: data = 8'hfe;
      17'd72177: data = 8'hfd;
      17'd72178: data = 8'hfe;
      17'd72179: data = 8'h01;
      17'd72180: data = 8'h00;
      17'd72181: data = 8'hfe;
      17'd72182: data = 8'hfe;
      17'd72183: data = 8'hfd;
      17'd72184: data = 8'hfe;
      17'd72185: data = 8'hfc;
      17'd72186: data = 8'hfc;
      17'd72187: data = 8'hfe;
      17'd72188: data = 8'hfd;
      17'd72189: data = 8'hfe;
      17'd72190: data = 8'hfd;
      17'd72191: data = 8'hfe;
      17'd72192: data = 8'h00;
      17'd72193: data = 8'h00;
      17'd72194: data = 8'h00;
      17'd72195: data = 8'h00;
      17'd72196: data = 8'h00;
      17'd72197: data = 8'h00;
      17'd72198: data = 8'hfe;
      17'd72199: data = 8'hfe;
      17'd72200: data = 8'hfe;
      17'd72201: data = 8'hfe;
      17'd72202: data = 8'hfe;
      17'd72203: data = 8'hfe;
      17'd72204: data = 8'h00;
      17'd72205: data = 8'h01;
      17'd72206: data = 8'h01;
      17'd72207: data = 8'h01;
      17'd72208: data = 8'h01;
      17'd72209: data = 8'h01;
      17'd72210: data = 8'h02;
      17'd72211: data = 8'h00;
      17'd72212: data = 8'hfe;
      17'd72213: data = 8'hfe;
      17'd72214: data = 8'hfd;
      17'd72215: data = 8'h00;
      17'd72216: data = 8'h00;
      17'd72217: data = 8'h01;
      17'd72218: data = 8'h01;
      17'd72219: data = 8'h01;
      17'd72220: data = 8'h04;
      17'd72221: data = 8'h05;
      17'd72222: data = 8'h04;
      17'd72223: data = 8'h04;
      17'd72224: data = 8'h04;
      17'd72225: data = 8'h02;
      17'd72226: data = 8'h02;
      17'd72227: data = 8'h01;
      17'd72228: data = 8'h00;
      17'd72229: data = 8'h00;
      17'd72230: data = 8'h00;
      17'd72231: data = 8'h01;
      17'd72232: data = 8'h00;
      17'd72233: data = 8'h00;
      17'd72234: data = 8'h00;
      17'd72235: data = 8'h00;
      17'd72236: data = 8'h00;
      17'd72237: data = 8'h00;
      17'd72238: data = 8'hfe;
      17'd72239: data = 8'hfd;
      17'd72240: data = 8'hfd;
      17'd72241: data = 8'hfd;
      17'd72242: data = 8'hfd;
      17'd72243: data = 8'hfc;
      17'd72244: data = 8'hfc;
      17'd72245: data = 8'hfd;
      17'd72246: data = 8'hfe;
      17'd72247: data = 8'hfe;
      17'd72248: data = 8'hfd;
      17'd72249: data = 8'hfe;
      17'd72250: data = 8'h00;
      17'd72251: data = 8'h01;
      17'd72252: data = 8'h01;
      17'd72253: data = 8'h00;
      17'd72254: data = 8'h00;
      17'd72255: data = 8'h00;
      17'd72256: data = 8'hfe;
      17'd72257: data = 8'hfe;
      17'd72258: data = 8'h01;
      17'd72259: data = 8'h00;
      17'd72260: data = 8'h00;
      17'd72261: data = 8'h01;
      17'd72262: data = 8'h01;
      17'd72263: data = 8'h00;
      17'd72264: data = 8'h01;
      17'd72265: data = 8'h02;
      17'd72266: data = 8'h04;
      17'd72267: data = 8'h05;
      17'd72268: data = 8'h05;
      17'd72269: data = 8'h02;
      17'd72270: data = 8'h02;
      17'd72271: data = 8'h04;
      17'd72272: data = 8'h01;
      17'd72273: data = 8'h01;
      17'd72274: data = 8'h01;
      17'd72275: data = 8'h01;
      17'd72276: data = 8'h01;
      17'd72277: data = 8'h01;
      17'd72278: data = 8'h00;
      17'd72279: data = 8'h01;
      17'd72280: data = 8'h02;
      17'd72281: data = 8'h01;
      17'd72282: data = 8'h02;
      17'd72283: data = 8'h02;
      17'd72284: data = 8'h02;
      17'd72285: data = 8'h00;
      17'd72286: data = 8'h00;
      17'd72287: data = 8'h01;
      17'd72288: data = 8'h00;
      17'd72289: data = 8'hfe;
      17'd72290: data = 8'h00;
      17'd72291: data = 8'h00;
      17'd72292: data = 8'h00;
      17'd72293: data = 8'h00;
      17'd72294: data = 8'h01;
      17'd72295: data = 8'h01;
      17'd72296: data = 8'h01;
      17'd72297: data = 8'h01;
      17'd72298: data = 8'hfe;
      17'd72299: data = 8'h01;
      17'd72300: data = 8'h00;
      17'd72301: data = 8'h00;
      17'd72302: data = 8'h00;
      17'd72303: data = 8'h00;
      17'd72304: data = 8'h00;
      17'd72305: data = 8'hfe;
      17'd72306: data = 8'h00;
      17'd72307: data = 8'h00;
      17'd72308: data = 8'hfe;
      17'd72309: data = 8'h00;
      17'd72310: data = 8'h00;
      17'd72311: data = 8'h00;
      17'd72312: data = 8'hfe;
      17'd72313: data = 8'hfd;
      17'd72314: data = 8'h00;
      17'd72315: data = 8'hfe;
      17'd72316: data = 8'hfc;
      17'd72317: data = 8'hfd;
      17'd72318: data = 8'hfd;
      17'd72319: data = 8'hfc;
      17'd72320: data = 8'hfe;
      17'd72321: data = 8'hfe;
      17'd72322: data = 8'hfe;
      17'd72323: data = 8'h00;
      17'd72324: data = 8'h01;
      17'd72325: data = 8'h01;
      17'd72326: data = 8'h00;
      17'd72327: data = 8'h01;
      17'd72328: data = 8'hfe;
      17'd72329: data = 8'hfe;
      17'd72330: data = 8'hfe;
      17'd72331: data = 8'hfe;
      17'd72332: data = 8'hfd;
      17'd72333: data = 8'hfd;
      17'd72334: data = 8'hfd;
      17'd72335: data = 8'hfe;
      17'd72336: data = 8'h00;
      17'd72337: data = 8'h00;
      17'd72338: data = 8'h01;
      17'd72339: data = 8'h01;
      17'd72340: data = 8'h01;
      17'd72341: data = 8'h01;
      17'd72342: data = 8'h02;
      17'd72343: data = 8'h02;
      17'd72344: data = 8'h01;
      17'd72345: data = 8'h00;
      17'd72346: data = 8'h00;
      17'd72347: data = 8'hfe;
      17'd72348: data = 8'h00;
      17'd72349: data = 8'h00;
      17'd72350: data = 8'hfe;
      17'd72351: data = 8'hfe;
      17'd72352: data = 8'hfe;
      17'd72353: data = 8'hfe;
      17'd72354: data = 8'h00;
      17'd72355: data = 8'h00;
      17'd72356: data = 8'h00;
      17'd72357: data = 8'h01;
      17'd72358: data = 8'h00;
      17'd72359: data = 8'h00;
      17'd72360: data = 8'hfe;
      17'd72361: data = 8'hfd;
      17'd72362: data = 8'hfd;
      17'd72363: data = 8'hfc;
      17'd72364: data = 8'hfc;
      17'd72365: data = 8'hfa;
      17'd72366: data = 8'hfc;
      17'd72367: data = 8'hfc;
      17'd72368: data = 8'hfa;
      17'd72369: data = 8'hfc;
      17'd72370: data = 8'hfd;
      17'd72371: data = 8'hfd;
      17'd72372: data = 8'hfe;
      17'd72373: data = 8'hfe;
      17'd72374: data = 8'hfd;
      17'd72375: data = 8'hfd;
      17'd72376: data = 8'hfd;
      17'd72377: data = 8'hfc;
      17'd72378: data = 8'hfd;
      17'd72379: data = 8'hfc;
      17'd72380: data = 8'hfa;
      17'd72381: data = 8'hfc;
      17'd72382: data = 8'hfc;
      17'd72383: data = 8'hfd;
      17'd72384: data = 8'hfe;
      17'd72385: data = 8'h00;
      17'd72386: data = 8'hfe;
      17'd72387: data = 8'h01;
      17'd72388: data = 8'h04;
      17'd72389: data = 8'h02;
      17'd72390: data = 8'h01;
      17'd72391: data = 8'h00;
      17'd72392: data = 8'h01;
      17'd72393: data = 8'h00;
      17'd72394: data = 8'hfe;
      17'd72395: data = 8'hfe;
      17'd72396: data = 8'hfc;
      17'd72397: data = 8'hfd;
      17'd72398: data = 8'hfc;
      17'd72399: data = 8'hfe;
      17'd72400: data = 8'h00;
      17'd72401: data = 8'h01;
      17'd72402: data = 8'h01;
      17'd72403: data = 8'h01;
      17'd72404: data = 8'h02;
      17'd72405: data = 8'h02;
      17'd72406: data = 8'h00;
      17'd72407: data = 8'hfe;
      17'd72408: data = 8'hfe;
      17'd72409: data = 8'hfe;
      17'd72410: data = 8'hfc;
      17'd72411: data = 8'hfc;
      17'd72412: data = 8'hfd;
      17'd72413: data = 8'hfd;
      17'd72414: data = 8'hfc;
      17'd72415: data = 8'hfd;
      17'd72416: data = 8'hfd;
      17'd72417: data = 8'hfc;
      17'd72418: data = 8'hfe;
      17'd72419: data = 8'hfd;
      17'd72420: data = 8'hfc;
      17'd72421: data = 8'hfe;
      17'd72422: data = 8'hfe;
      17'd72423: data = 8'hfc;
      17'd72424: data = 8'hfc;
      17'd72425: data = 8'hfc;
      17'd72426: data = 8'hfc;
      17'd72427: data = 8'hfa;
      17'd72428: data = 8'hfc;
      17'd72429: data = 8'hfd;
      17'd72430: data = 8'hfc;
      17'd72431: data = 8'hfd;
      17'd72432: data = 8'hfd;
      17'd72433: data = 8'hfd;
      17'd72434: data = 8'hfe;
      17'd72435: data = 8'hfd;
      17'd72436: data = 8'hfd;
      17'd72437: data = 8'hfd;
      17'd72438: data = 8'hfc;
      17'd72439: data = 8'hfc;
      17'd72440: data = 8'hfa;
      17'd72441: data = 8'hfa;
      17'd72442: data = 8'hfd;
      17'd72443: data = 8'hfc;
      17'd72444: data = 8'hfd;
      17'd72445: data = 8'hfc;
      17'd72446: data = 8'hfc;
      17'd72447: data = 8'hfd;
      17'd72448: data = 8'h00;
      17'd72449: data = 8'h00;
      17'd72450: data = 8'hfe;
      17'd72451: data = 8'h01;
      17'd72452: data = 8'hfe;
      17'd72453: data = 8'hfe;
      17'd72454: data = 8'h00;
      17'd72455: data = 8'hfe;
      17'd72456: data = 8'hfd;
      17'd72457: data = 8'hfd;
      17'd72458: data = 8'hfe;
      17'd72459: data = 8'hfe;
      17'd72460: data = 8'h00;
      17'd72461: data = 8'h00;
      17'd72462: data = 8'h00;
      17'd72463: data = 8'h01;
      17'd72464: data = 8'h02;
      17'd72465: data = 8'h04;
      17'd72466: data = 8'h02;
      17'd72467: data = 8'h01;
      17'd72468: data = 8'h01;
      17'd72469: data = 8'h04;
      17'd72470: data = 8'h02;
      17'd72471: data = 8'h01;
      17'd72472: data = 8'h00;
      17'd72473: data = 8'h01;
      17'd72474: data = 8'h00;
      17'd72475: data = 8'h00;
      17'd72476: data = 8'h00;
      17'd72477: data = 8'hfe;
      17'd72478: data = 8'h01;
      17'd72479: data = 8'h02;
      17'd72480: data = 8'h01;
      17'd72481: data = 8'h01;
      17'd72482: data = 8'h01;
      17'd72483: data = 8'h00;
      17'd72484: data = 8'h00;
      17'd72485: data = 8'hfe;
      17'd72486: data = 8'hfe;
      17'd72487: data = 8'hfc;
      17'd72488: data = 8'hfc;
      17'd72489: data = 8'hfd;
      17'd72490: data = 8'hfc;
      17'd72491: data = 8'hfd;
      17'd72492: data = 8'hfd;
      17'd72493: data = 8'hfe;
      17'd72494: data = 8'h00;
      17'd72495: data = 8'h00;
      17'd72496: data = 8'hfe;
      17'd72497: data = 8'h00;
      17'd72498: data = 8'h00;
      17'd72499: data = 8'hfe;
      17'd72500: data = 8'h01;
      17'd72501: data = 8'hfe;
      17'd72502: data = 8'hfe;
      17'd72503: data = 8'h00;
      17'd72504: data = 8'hfe;
      17'd72505: data = 8'hfe;
      17'd72506: data = 8'h00;
      17'd72507: data = 8'hfe;
      17'd72508: data = 8'h00;
      17'd72509: data = 8'h00;
      17'd72510: data = 8'h01;
      17'd72511: data = 8'h02;
      17'd72512: data = 8'h02;
      17'd72513: data = 8'h02;
      17'd72514: data = 8'h02;
      17'd72515: data = 8'h04;
      17'd72516: data = 8'h02;
      17'd72517: data = 8'h04;
      17'd72518: data = 8'h02;
      17'd72519: data = 8'h01;
      17'd72520: data = 8'hfe;
      17'd72521: data = 8'h01;
      17'd72522: data = 8'h01;
      17'd72523: data = 8'h01;
      17'd72524: data = 8'h02;
      17'd72525: data = 8'h02;
      17'd72526: data = 8'h02;
      17'd72527: data = 8'h01;
      17'd72528: data = 8'h01;
      17'd72529: data = 8'h00;
      17'd72530: data = 8'h01;
      17'd72531: data = 8'h01;
      17'd72532: data = 8'h00;
      17'd72533: data = 8'h00;
      17'd72534: data = 8'h01;
      17'd72535: data = 8'hfe;
      17'd72536: data = 8'hfe;
      17'd72537: data = 8'hfe;
      17'd72538: data = 8'hfe;
      17'd72539: data = 8'hfe;
      17'd72540: data = 8'hfe;
      17'd72541: data = 8'h00;
      17'd72542: data = 8'h01;
      17'd72543: data = 8'h01;
      17'd72544: data = 8'h02;
      17'd72545: data = 8'h01;
      17'd72546: data = 8'h00;
      17'd72547: data = 8'h01;
      17'd72548: data = 8'h01;
      17'd72549: data = 8'h01;
      17'd72550: data = 8'h00;
      17'd72551: data = 8'hfe;
      17'd72552: data = 8'h01;
      17'd72553: data = 8'h00;
      17'd72554: data = 8'hfd;
      17'd72555: data = 8'h00;
      17'd72556: data = 8'h00;
      17'd72557: data = 8'h00;
      17'd72558: data = 8'h01;
      17'd72559: data = 8'hfe;
      17'd72560: data = 8'hfe;
      17'd72561: data = 8'h00;
      17'd72562: data = 8'h00;
      17'd72563: data = 8'h00;
      17'd72564: data = 8'h01;
      17'd72565: data = 8'h02;
      17'd72566: data = 8'h02;
      17'd72567: data = 8'h01;
      17'd72568: data = 8'h01;
      17'd72569: data = 8'h01;
      17'd72570: data = 8'h01;
      17'd72571: data = 8'h01;
      17'd72572: data = 8'hfe;
      17'd72573: data = 8'h00;
      17'd72574: data = 8'h00;
      17'd72575: data = 8'hfe;
      17'd72576: data = 8'hfe;
      17'd72577: data = 8'h00;
      17'd72578: data = 8'h00;
      17'd72579: data = 8'h00;
      17'd72580: data = 8'h00;
      17'd72581: data = 8'h00;
      17'd72582: data = 8'hfe;
      17'd72583: data = 8'hfe;
      17'd72584: data = 8'hfe;
      17'd72585: data = 8'hfd;
      17'd72586: data = 8'h00;
      17'd72587: data = 8'h01;
      17'd72588: data = 8'h00;
      17'd72589: data = 8'h00;
      17'd72590: data = 8'hfd;
      17'd72591: data = 8'hfc;
      17'd72592: data = 8'hfe;
      17'd72593: data = 8'hfe;
      17'd72594: data = 8'hfe;
      17'd72595: data = 8'hfe;
      17'd72596: data = 8'hfe;
      17'd72597: data = 8'hfe;
      17'd72598: data = 8'hfd;
      17'd72599: data = 8'hfe;
      17'd72600: data = 8'hfd;
      17'd72601: data = 8'hfe;
      17'd72602: data = 8'h00;
      17'd72603: data = 8'h00;
      17'd72604: data = 8'h00;
      17'd72605: data = 8'hfe;
      17'd72606: data = 8'hfe;
      17'd72607: data = 8'h00;
      17'd72608: data = 8'hfe;
      17'd72609: data = 8'hfe;
      17'd72610: data = 8'h00;
      17'd72611: data = 8'hfe;
      17'd72612: data = 8'h00;
      17'd72613: data = 8'h02;
      17'd72614: data = 8'h00;
      17'd72615: data = 8'h00;
      17'd72616: data = 8'h02;
      17'd72617: data = 8'h02;
      17'd72618: data = 8'h01;
      17'd72619: data = 8'h00;
      17'd72620: data = 8'hfe;
      17'd72621: data = 8'hfe;
      17'd72622: data = 8'hfe;
      17'd72623: data = 8'hfe;
      17'd72624: data = 8'h00;
      17'd72625: data = 8'h01;
      17'd72626: data = 8'h01;
      17'd72627: data = 8'hfe;
      17'd72628: data = 8'hfe;
      17'd72629: data = 8'hfe;
      17'd72630: data = 8'hfe;
      17'd72631: data = 8'hfe;
      17'd72632: data = 8'hfe;
      17'd72633: data = 8'h00;
      17'd72634: data = 8'hfe;
      17'd72635: data = 8'hfe;
      17'd72636: data = 8'hfe;
      17'd72637: data = 8'hfd;
      17'd72638: data = 8'hfd;
      17'd72639: data = 8'hfd;
      17'd72640: data = 8'hfe;
      17'd72641: data = 8'hfe;
      17'd72642: data = 8'hfe;
      17'd72643: data = 8'hfe;
      17'd72644: data = 8'h00;
      17'd72645: data = 8'h00;
      17'd72646: data = 8'h00;
      17'd72647: data = 8'h00;
      17'd72648: data = 8'h00;
      17'd72649: data = 8'h00;
      17'd72650: data = 8'h01;
      17'd72651: data = 8'h00;
      17'd72652: data = 8'h00;
      17'd72653: data = 8'h04;
      17'd72654: data = 8'h02;
      17'd72655: data = 8'h02;
      17'd72656: data = 8'h04;
      17'd72657: data = 8'h02;
      17'd72658: data = 8'h02;
      17'd72659: data = 8'h01;
      17'd72660: data = 8'h01;
      17'd72661: data = 8'h00;
      17'd72662: data = 8'h00;
      17'd72663: data = 8'h01;
      17'd72664: data = 8'h00;
      17'd72665: data = 8'h04;
      17'd72666: data = 8'h01;
      17'd72667: data = 8'h01;
      17'd72668: data = 8'h01;
      17'd72669: data = 8'h00;
      17'd72670: data = 8'h01;
      17'd72671: data = 8'h00;
      17'd72672: data = 8'hfe;
      17'd72673: data = 8'hfd;
      17'd72674: data = 8'hfd;
      17'd72675: data = 8'hfa;
      17'd72676: data = 8'hfd;
      17'd72677: data = 8'hfd;
      17'd72678: data = 8'hfd;
      17'd72679: data = 8'hfd;
      17'd72680: data = 8'hfd;
      17'd72681: data = 8'hfd;
      17'd72682: data = 8'hfd;
      17'd72683: data = 8'hfd;
      17'd72684: data = 8'hfc;
      17'd72685: data = 8'hfc;
      17'd72686: data = 8'hfe;
      17'd72687: data = 8'hfd;
      17'd72688: data = 8'hfd;
      17'd72689: data = 8'hfd;
      17'd72690: data = 8'hfd;
      17'd72691: data = 8'hfd;
      17'd72692: data = 8'hfd;
      17'd72693: data = 8'hfe;
      17'd72694: data = 8'hfc;
      17'd72695: data = 8'hfe;
      17'd72696: data = 8'h00;
      17'd72697: data = 8'h00;
      17'd72698: data = 8'hfe;
      17'd72699: data = 8'hfe;
      17'd72700: data = 8'hfe;
      17'd72701: data = 8'hfe;
      17'd72702: data = 8'h01;
      17'd72703: data = 8'h00;
      17'd72704: data = 8'h01;
      17'd72705: data = 8'h01;
      17'd72706: data = 8'h01;
      17'd72707: data = 8'h02;
      17'd72708: data = 8'h02;
      17'd72709: data = 8'h01;
      17'd72710: data = 8'h00;
      17'd72711: data = 8'h00;
      17'd72712: data = 8'h00;
      17'd72713: data = 8'h02;
      17'd72714: data = 8'h01;
      17'd72715: data = 8'h01;
      17'd72716: data = 8'h02;
      17'd72717: data = 8'h02;
      17'd72718: data = 8'h01;
      17'd72719: data = 8'h01;
      17'd72720: data = 8'h01;
      17'd72721: data = 8'h00;
      17'd72722: data = 8'h01;
      17'd72723: data = 8'h00;
      17'd72724: data = 8'h00;
      17'd72725: data = 8'h00;
      17'd72726: data = 8'hfe;
      17'd72727: data = 8'hfe;
      17'd72728: data = 8'hfe;
      17'd72729: data = 8'h00;
      17'd72730: data = 8'hfe;
      17'd72731: data = 8'hfe;
      17'd72732: data = 8'h00;
      17'd72733: data = 8'h00;
      17'd72734: data = 8'hfe;
      17'd72735: data = 8'hfd;
      17'd72736: data = 8'hfe;
      17'd72737: data = 8'hfd;
      17'd72738: data = 8'hfd;
      17'd72739: data = 8'hfe;
      17'd72740: data = 8'hfd;
      17'd72741: data = 8'hfd;
      17'd72742: data = 8'hfe;
      17'd72743: data = 8'h00;
      17'd72744: data = 8'h00;
      17'd72745: data = 8'hfe;
      17'd72746: data = 8'h01;
      17'd72747: data = 8'h00;
      17'd72748: data = 8'hfe;
      17'd72749: data = 8'hfe;
      17'd72750: data = 8'hfe;
      17'd72751: data = 8'h00;
      17'd72752: data = 8'hfe;
      17'd72753: data = 8'h01;
      17'd72754: data = 8'h01;
      17'd72755: data = 8'h00;
      17'd72756: data = 8'h00;
      17'd72757: data = 8'h00;
      17'd72758: data = 8'h02;
      17'd72759: data = 8'h01;
      17'd72760: data = 8'h00;
      17'd72761: data = 8'hfe;
      17'd72762: data = 8'hfe;
      17'd72763: data = 8'h00;
      17'd72764: data = 8'h00;
      17'd72765: data = 8'hfe;
      17'd72766: data = 8'h00;
      17'd72767: data = 8'hfe;
      17'd72768: data = 8'hfe;
      17'd72769: data = 8'hfd;
      17'd72770: data = 8'hfe;
      17'd72771: data = 8'hfe;
      17'd72772: data = 8'hfe;
      17'd72773: data = 8'h00;
      17'd72774: data = 8'h00;
      17'd72775: data = 8'h00;
      17'd72776: data = 8'hfe;
      17'd72777: data = 8'h00;
      17'd72778: data = 8'h00;
      17'd72779: data = 8'h00;
      17'd72780: data = 8'h00;
      17'd72781: data = 8'hfe;
      17'd72782: data = 8'hfd;
      17'd72783: data = 8'hfe;
      17'd72784: data = 8'hfe;
      17'd72785: data = 8'hfd;
      17'd72786: data = 8'hfe;
      17'd72787: data = 8'h00;
      17'd72788: data = 8'hfe;
      17'd72789: data = 8'hfe;
      17'd72790: data = 8'h00;
      17'd72791: data = 8'hfe;
      17'd72792: data = 8'h00;
      17'd72793: data = 8'h01;
      17'd72794: data = 8'h00;
      17'd72795: data = 8'hfe;
      17'd72796: data = 8'hfe;
      17'd72797: data = 8'hfd;
      17'd72798: data = 8'hfd;
      17'd72799: data = 8'hfc;
      17'd72800: data = 8'hfd;
      17'd72801: data = 8'hfd;
      17'd72802: data = 8'hfd;
      17'd72803: data = 8'hfe;
      17'd72804: data = 8'hfe;
      17'd72805: data = 8'hfe;
      17'd72806: data = 8'h00;
      17'd72807: data = 8'h00;
      17'd72808: data = 8'hfe;
      17'd72809: data = 8'hfd;
      17'd72810: data = 8'hfe;
      17'd72811: data = 8'hfd;
      17'd72812: data = 8'hfd;
      17'd72813: data = 8'hfe;
      17'd72814: data = 8'hfe;
      17'd72815: data = 8'h00;
      17'd72816: data = 8'h00;
      17'd72817: data = 8'h01;
      17'd72818: data = 8'h01;
      17'd72819: data = 8'h01;
      17'd72820: data = 8'h01;
      17'd72821: data = 8'h01;
      17'd72822: data = 8'h01;
      17'd72823: data = 8'h02;
      17'd72824: data = 8'h02;
      17'd72825: data = 8'h01;
      17'd72826: data = 8'h02;
      17'd72827: data = 8'h02;
      17'd72828: data = 8'h04;
      17'd72829: data = 8'h04;
      17'd72830: data = 8'h02;
      17'd72831: data = 8'h04;
      17'd72832: data = 8'h02;
      17'd72833: data = 8'h02;
      17'd72834: data = 8'h01;
      17'd72835: data = 8'h04;
      17'd72836: data = 8'h01;
      17'd72837: data = 8'h00;
      17'd72838: data = 8'h00;
      17'd72839: data = 8'h00;
      17'd72840: data = 8'h00;
      17'd72841: data = 8'h01;
      17'd72842: data = 8'h00;
      17'd72843: data = 8'h00;
      17'd72844: data = 8'h00;
      17'd72845: data = 8'hfe;
      17'd72846: data = 8'h00;
      17'd72847: data = 8'h01;
      17'd72848: data = 8'h00;
      17'd72849: data = 8'h00;
      17'd72850: data = 8'hfe;
      17'd72851: data = 8'hfe;
      17'd72852: data = 8'hfe;
      17'd72853: data = 8'hfd;
      17'd72854: data = 8'hfd;
      17'd72855: data = 8'hfa;
      17'd72856: data = 8'hfa;
      17'd72857: data = 8'hfd;
      17'd72858: data = 8'hfd;
      17'd72859: data = 8'hfc;
      17'd72860: data = 8'hfd;
      17'd72861: data = 8'hfd;
      17'd72862: data = 8'hfc;
      17'd72863: data = 8'hfd;
      17'd72864: data = 8'hfd;
      17'd72865: data = 8'hfe;
      17'd72866: data = 8'h00;
      17'd72867: data = 8'h00;
      17'd72868: data = 8'hfe;
      17'd72869: data = 8'h00;
      17'd72870: data = 8'hfe;
      17'd72871: data = 8'hfe;
      17'd72872: data = 8'h00;
      17'd72873: data = 8'hfe;
      17'd72874: data = 8'hfe;
      17'd72875: data = 8'hfe;
      17'd72876: data = 8'hfe;
      17'd72877: data = 8'h00;
      17'd72878: data = 8'h00;
      17'd72879: data = 8'h00;
      17'd72880: data = 8'h00;
      17'd72881: data = 8'h00;
      17'd72882: data = 8'h01;
      17'd72883: data = 8'h01;
      17'd72884: data = 8'h04;
      17'd72885: data = 8'h02;
      17'd72886: data = 8'h00;
      17'd72887: data = 8'h01;
      17'd72888: data = 8'h00;
      17'd72889: data = 8'hfe;
      17'd72890: data = 8'h00;
      17'd72891: data = 8'h01;
      17'd72892: data = 8'h00;
      17'd72893: data = 8'h01;
      17'd72894: data = 8'h02;
      17'd72895: data = 8'h02;
      17'd72896: data = 8'h02;
      17'd72897: data = 8'h02;
      17'd72898: data = 8'h01;
      17'd72899: data = 8'h00;
      17'd72900: data = 8'h00;
      17'd72901: data = 8'h01;
      17'd72902: data = 8'h00;
      17'd72903: data = 8'h01;
      17'd72904: data = 8'h00;
      17'd72905: data = 8'hfe;
      17'd72906: data = 8'hfc;
      17'd72907: data = 8'hfa;
      17'd72908: data = 8'hfd;
      17'd72909: data = 8'hfd;
      17'd72910: data = 8'hfc;
      17'd72911: data = 8'hfe;
      17'd72912: data = 8'hfe;
      17'd72913: data = 8'hfe;
      17'd72914: data = 8'hfd;
      17'd72915: data = 8'hfd;
      17'd72916: data = 8'hfc;
      17'd72917: data = 8'hfa;
      17'd72918: data = 8'hfc;
      17'd72919: data = 8'hfa;
      17'd72920: data = 8'hfa;
      17'd72921: data = 8'hfc;
      17'd72922: data = 8'hfd;
      17'd72923: data = 8'hfc;
      17'd72924: data = 8'hfd;
      17'd72925: data = 8'hfe;
      17'd72926: data = 8'hfd;
      17'd72927: data = 8'hfd;
      17'd72928: data = 8'hfd;
      17'd72929: data = 8'hfd;
      17'd72930: data = 8'h01;
      17'd72931: data = 8'h01;
      17'd72932: data = 8'h00;
      17'd72933: data = 8'h00;
      17'd72934: data = 8'hfe;
      17'd72935: data = 8'hfe;
      17'd72936: data = 8'h00;
      17'd72937: data = 8'hfe;
      17'd72938: data = 8'hfd;
      17'd72939: data = 8'hfe;
      17'd72940: data = 8'hfe;
      17'd72941: data = 8'hfe;
      17'd72942: data = 8'h00;
      17'd72943: data = 8'h00;
      17'd72944: data = 8'h00;
      17'd72945: data = 8'h01;
      17'd72946: data = 8'h01;
      17'd72947: data = 8'h00;
      17'd72948: data = 8'h01;
      17'd72949: data = 8'h01;
      17'd72950: data = 8'hfe;
      17'd72951: data = 8'hfe;
      17'd72952: data = 8'hfe;
      17'd72953: data = 8'hfd;
      17'd72954: data = 8'h00;
      17'd72955: data = 8'h00;
      17'd72956: data = 8'hfe;
      17'd72957: data = 8'h00;
      17'd72958: data = 8'h02;
      17'd72959: data = 8'h00;
      17'd72960: data = 8'h00;
      17'd72961: data = 8'h01;
      17'd72962: data = 8'h00;
      17'd72963: data = 8'hfe;
      17'd72964: data = 8'hfd;
      17'd72965: data = 8'hfe;
      17'd72966: data = 8'hfe;
      17'd72967: data = 8'hfd;
      17'd72968: data = 8'hfd;
      17'd72969: data = 8'h00;
      17'd72970: data = 8'hfe;
      17'd72971: data = 8'h00;
      17'd72972: data = 8'h00;
      17'd72973: data = 8'h00;
      17'd72974: data = 8'h00;
      17'd72975: data = 8'h00;
      17'd72976: data = 8'h01;
      17'd72977: data = 8'hfd;
      17'd72978: data = 8'hfe;
      17'd72979: data = 8'h00;
      17'd72980: data = 8'hfe;
      17'd72981: data = 8'hfe;
      17'd72982: data = 8'h01;
      17'd72983: data = 8'h01;
      17'd72984: data = 8'h01;
      17'd72985: data = 8'h00;
      17'd72986: data = 8'h00;
      17'd72987: data = 8'h01;
      17'd72988: data = 8'h01;
      17'd72989: data = 8'h01;
      17'd72990: data = 8'h01;
      17'd72991: data = 8'h01;
      17'd72992: data = 8'h02;
      17'd72993: data = 8'h01;
      17'd72994: data = 8'hfe;
      17'd72995: data = 8'h00;
      17'd72996: data = 8'h00;
      17'd72997: data = 8'h01;
      17'd72998: data = 8'h01;
      17'd72999: data = 8'h01;
      17'd73000: data = 8'h02;
      17'd73001: data = 8'h01;
      17'd73002: data = 8'h01;
      17'd73003: data = 8'h01;
      17'd73004: data = 8'h00;
      17'd73005: data = 8'h00;
      17'd73006: data = 8'h00;
      17'd73007: data = 8'h01;
      17'd73008: data = 8'h00;
      17'd73009: data = 8'h00;
      17'd73010: data = 8'h01;
      17'd73011: data = 8'h00;
      17'd73012: data = 8'h01;
      17'd73013: data = 8'h02;
      17'd73014: data = 8'h01;
      17'd73015: data = 8'h01;
      17'd73016: data = 8'h02;
      17'd73017: data = 8'h01;
      17'd73018: data = 8'h02;
      17'd73019: data = 8'h01;
      17'd73020: data = 8'h00;
      17'd73021: data = 8'hfe;
      17'd73022: data = 8'h00;
      17'd73023: data = 8'h00;
      17'd73024: data = 8'hfe;
      17'd73025: data = 8'h01;
      17'd73026: data = 8'hfe;
      17'd73027: data = 8'hfe;
      17'd73028: data = 8'h00;
      17'd73029: data = 8'h00;
      17'd73030: data = 8'h01;
      17'd73031: data = 8'h00;
      17'd73032: data = 8'h00;
      17'd73033: data = 8'hfe;
      17'd73034: data = 8'hfe;
      17'd73035: data = 8'h00;
      17'd73036: data = 8'h00;
      17'd73037: data = 8'h00;
      17'd73038: data = 8'hfe;
      17'd73039: data = 8'h00;
      17'd73040: data = 8'h01;
      17'd73041: data = 8'h00;
      17'd73042: data = 8'h00;
      17'd73043: data = 8'h01;
      17'd73044: data = 8'h01;
      17'd73045: data = 8'h01;
      17'd73046: data = 8'h01;
      17'd73047: data = 8'h00;
      17'd73048: data = 8'hfe;
      17'd73049: data = 8'hfe;
      17'd73050: data = 8'h00;
      17'd73051: data = 8'hfe;
      17'd73052: data = 8'h01;
      17'd73053: data = 8'hfe;
      17'd73054: data = 8'hfe;
      17'd73055: data = 8'h00;
      17'd73056: data = 8'hfe;
      17'd73057: data = 8'h01;
      17'd73058: data = 8'h01;
      17'd73059: data = 8'h02;
      17'd73060: data = 8'h01;
      17'd73061: data = 8'h01;
      17'd73062: data = 8'h02;
      17'd73063: data = 8'h00;
      17'd73064: data = 8'h01;
      17'd73065: data = 8'h00;
      17'd73066: data = 8'hfd;
      17'd73067: data = 8'hfd;
      17'd73068: data = 8'hfe;
      17'd73069: data = 8'hfe;
      17'd73070: data = 8'h00;
      17'd73071: data = 8'h00;
      17'd73072: data = 8'h01;
      17'd73073: data = 8'h01;
      17'd73074: data = 8'h02;
      17'd73075: data = 8'h01;
      17'd73076: data = 8'h01;
      17'd73077: data = 8'h01;
      17'd73078: data = 8'h00;
      17'd73079: data = 8'h01;
      17'd73080: data = 8'h01;
      17'd73081: data = 8'h00;
      17'd73082: data = 8'h00;
      17'd73083: data = 8'h00;
      17'd73084: data = 8'h00;
      17'd73085: data = 8'h01;
      17'd73086: data = 8'h02;
      17'd73087: data = 8'h01;
      17'd73088: data = 8'h01;
      17'd73089: data = 8'h04;
      17'd73090: data = 8'h01;
      17'd73091: data = 8'h01;
      17'd73092: data = 8'h02;
      17'd73093: data = 8'h00;
      17'd73094: data = 8'h00;
      17'd73095: data = 8'hfd;
      17'd73096: data = 8'hfd;
      17'd73097: data = 8'hfe;
      17'd73098: data = 8'hfe;
      17'd73099: data = 8'hfd;
      17'd73100: data = 8'h00;
      17'd73101: data = 8'h02;
      17'd73102: data = 8'h00;
      17'd73103: data = 8'h01;
      17'd73104: data = 8'h02;
      17'd73105: data = 8'hfe;
      17'd73106: data = 8'h00;
      17'd73107: data = 8'h01;
      17'd73108: data = 8'hfd;
      17'd73109: data = 8'h00;
      17'd73110: data = 8'hfe;
      17'd73111: data = 8'hfd;
      17'd73112: data = 8'hfe;
      17'd73113: data = 8'hfd;
      17'd73114: data = 8'hfe;
      17'd73115: data = 8'hfd;
      17'd73116: data = 8'hfe;
      17'd73117: data = 8'h01;
      17'd73118: data = 8'hfe;
      17'd73119: data = 8'h00;
      17'd73120: data = 8'h02;
      17'd73121: data = 8'h00;
      17'd73122: data = 8'h01;
      17'd73123: data = 8'h00;
      17'd73124: data = 8'hfd;
      17'd73125: data = 8'hfe;
      17'd73126: data = 8'h00;
      17'd73127: data = 8'hfd;
      17'd73128: data = 8'hfe;
      17'd73129: data = 8'h00;
      17'd73130: data = 8'h00;
      17'd73131: data = 8'h01;
      17'd73132: data = 8'h02;
      17'd73133: data = 8'h02;
      17'd73134: data = 8'h04;
      17'd73135: data = 8'h04;
      17'd73136: data = 8'h01;
      17'd73137: data = 8'h02;
      17'd73138: data = 8'h02;
      17'd73139: data = 8'h01;
      17'd73140: data = 8'h02;
      17'd73141: data = 8'h02;
      17'd73142: data = 8'h01;
      17'd73143: data = 8'h00;
      17'd73144: data = 8'h00;
      17'd73145: data = 8'hfe;
      17'd73146: data = 8'h00;
      17'd73147: data = 8'h01;
      17'd73148: data = 8'h00;
      17'd73149: data = 8'h00;
      17'd73150: data = 8'h01;
      17'd73151: data = 8'h00;
      17'd73152: data = 8'hfe;
      17'd73153: data = 8'h00;
      17'd73154: data = 8'hfe;
      17'd73155: data = 8'hfe;
      17'd73156: data = 8'h00;
      17'd73157: data = 8'hfd;
      17'd73158: data = 8'hfa;
      17'd73159: data = 8'hfa;
      17'd73160: data = 8'hfc;
      17'd73161: data = 8'hfd;
      17'd73162: data = 8'hfd;
      17'd73163: data = 8'hfd;
      17'd73164: data = 8'hfd;
      17'd73165: data = 8'hfd;
      17'd73166: data = 8'hfd;
      17'd73167: data = 8'hfd;
      17'd73168: data = 8'hfd;
      17'd73169: data = 8'hfd;
      17'd73170: data = 8'hfd;
      17'd73171: data = 8'hfe;
      17'd73172: data = 8'hfe;
      17'd73173: data = 8'hfe;
      17'd73174: data = 8'h00;
      17'd73175: data = 8'hfe;
      17'd73176: data = 8'hfd;
      17'd73177: data = 8'h02;
      17'd73178: data = 8'h01;
      17'd73179: data = 8'h00;
      17'd73180: data = 8'h01;
      17'd73181: data = 8'h01;
      17'd73182: data = 8'h01;
      17'd73183: data = 8'h00;
      17'd73184: data = 8'h00;
      17'd73185: data = 8'hfe;
      17'd73186: data = 8'hfe;
      17'd73187: data = 8'h01;
      17'd73188: data = 8'hfe;
      17'd73189: data = 8'hfd;
      17'd73190: data = 8'h01;
      17'd73191: data = 8'h01;
      17'd73192: data = 8'h01;
      17'd73193: data = 8'h02;
      17'd73194: data = 8'h00;
      17'd73195: data = 8'h00;
      17'd73196: data = 8'h01;
      17'd73197: data = 8'h00;
      17'd73198: data = 8'hfd;
      17'd73199: data = 8'hfc;
      17'd73200: data = 8'hfc;
      17'd73201: data = 8'hfc;
      17'd73202: data = 8'hfd;
      17'd73203: data = 8'hfe;
      17'd73204: data = 8'hfd;
      17'd73205: data = 8'h00;
      17'd73206: data = 8'h00;
      17'd73207: data = 8'h00;
      17'd73208: data = 8'h01;
      17'd73209: data = 8'hfe;
      17'd73210: data = 8'hfe;
      17'd73211: data = 8'h00;
      17'd73212: data = 8'hfd;
      17'd73213: data = 8'hfd;
      17'd73214: data = 8'hfd;
      17'd73215: data = 8'hfd;
      17'd73216: data = 8'hfd;
      17'd73217: data = 8'hfd;
      17'd73218: data = 8'hfe;
      17'd73219: data = 8'hfd;
      17'd73220: data = 8'h00;
      17'd73221: data = 8'h01;
      17'd73222: data = 8'h00;
      17'd73223: data = 8'h02;
      17'd73224: data = 8'h00;
      17'd73225: data = 8'h00;
      17'd73226: data = 8'h00;
      17'd73227: data = 8'h00;
      17'd73228: data = 8'hfe;
      17'd73229: data = 8'hfe;
      17'd73230: data = 8'hfe;
      17'd73231: data = 8'hfe;
      17'd73232: data = 8'hfe;
      17'd73233: data = 8'hfc;
      17'd73234: data = 8'hfc;
      17'd73235: data = 8'hfe;
      17'd73236: data = 8'h01;
      17'd73237: data = 8'h01;
      17'd73238: data = 8'h01;
      17'd73239: data = 8'h01;
      17'd73240: data = 8'h02;
      17'd73241: data = 8'h01;
      17'd73242: data = 8'h01;
      17'd73243: data = 8'h00;
      17'd73244: data = 8'hfd;
      17'd73245: data = 8'hfd;
      17'd73246: data = 8'hfd;
      17'd73247: data = 8'hfe;
      17'd73248: data = 8'h00;
      17'd73249: data = 8'h00;
      17'd73250: data = 8'h00;
      17'd73251: data = 8'h01;
      17'd73252: data = 8'h01;
      17'd73253: data = 8'h00;
      17'd73254: data = 8'h01;
      17'd73255: data = 8'h00;
      17'd73256: data = 8'h00;
      17'd73257: data = 8'h01;
      17'd73258: data = 8'hfe;
      17'd73259: data = 8'hfe;
      17'd73260: data = 8'h00;
      17'd73261: data = 8'hfe;
      17'd73262: data = 8'hfe;
      17'd73263: data = 8'hfe;
      17'd73264: data = 8'hfd;
      17'd73265: data = 8'h00;
      17'd73266: data = 8'h00;
      17'd73267: data = 8'hfe;
      17'd73268: data = 8'h00;
      17'd73269: data = 8'h00;
      17'd73270: data = 8'hfe;
      17'd73271: data = 8'hfd;
      17'd73272: data = 8'hfe;
      17'd73273: data = 8'hfd;
      17'd73274: data = 8'hfe;
      17'd73275: data = 8'hfd;
      17'd73276: data = 8'hfd;
      17'd73277: data = 8'hfe;
      17'd73278: data = 8'hfe;
      17'd73279: data = 8'hfd;
      17'd73280: data = 8'hfd;
      17'd73281: data = 8'h00;
      17'd73282: data = 8'h00;
      17'd73283: data = 8'hfd;
      17'd73284: data = 8'hfe;
      17'd73285: data = 8'hfd;
      17'd73286: data = 8'hfd;
      17'd73287: data = 8'h00;
      17'd73288: data = 8'hfe;
      17'd73289: data = 8'hfe;
      17'd73290: data = 8'hfd;
      17'd73291: data = 8'hfd;
      17'd73292: data = 8'hfd;
      17'd73293: data = 8'hfe;
      17'd73294: data = 8'h00;
      17'd73295: data = 8'h00;
      17'd73296: data = 8'h00;
      17'd73297: data = 8'h00;
      17'd73298: data = 8'h00;
      17'd73299: data = 8'h00;
      17'd73300: data = 8'h01;
      17'd73301: data = 8'h00;
      17'd73302: data = 8'h01;
      17'd73303: data = 8'h00;
      17'd73304: data = 8'hfe;
      17'd73305: data = 8'hfe;
      17'd73306: data = 8'hfe;
      17'd73307: data = 8'h00;
      17'd73308: data = 8'hfe;
      17'd73309: data = 8'h00;
      17'd73310: data = 8'h00;
      17'd73311: data = 8'h01;
      17'd73312: data = 8'h01;
      17'd73313: data = 8'h01;
      17'd73314: data = 8'h01;
      17'd73315: data = 8'h00;
      17'd73316: data = 8'h00;
      17'd73317: data = 8'hfe;
      17'd73318: data = 8'h00;
      17'd73319: data = 8'hfe;
      17'd73320: data = 8'hfd;
      17'd73321: data = 8'hfe;
      17'd73322: data = 8'h00;
      17'd73323: data = 8'hfd;
      17'd73324: data = 8'hfe;
      17'd73325: data = 8'hfe;
      17'd73326: data = 8'hfd;
      17'd73327: data = 8'h00;
      17'd73328: data = 8'hfe;
      17'd73329: data = 8'hfd;
      17'd73330: data = 8'hfe;
      17'd73331: data = 8'hfe;
      17'd73332: data = 8'hfe;
      17'd73333: data = 8'h00;
      17'd73334: data = 8'hfe;
      17'd73335: data = 8'hfd;
      17'd73336: data = 8'hfd;
      17'd73337: data = 8'hfd;
      17'd73338: data = 8'hfe;
      17'd73339: data = 8'hfd;
      17'd73340: data = 8'hfd;
      17'd73341: data = 8'hfd;
      17'd73342: data = 8'h00;
      17'd73343: data = 8'h00;
      17'd73344: data = 8'hfd;
      17'd73345: data = 8'h00;
      17'd73346: data = 8'h01;
      17'd73347: data = 8'h00;
      17'd73348: data = 8'h00;
      17'd73349: data = 8'h00;
      17'd73350: data = 8'hfe;
      17'd73351: data = 8'hfe;
      17'd73352: data = 8'hfe;
      17'd73353: data = 8'hfe;
      17'd73354: data = 8'hfe;
      17'd73355: data = 8'hfe;
      17'd73356: data = 8'hfe;
      17'd73357: data = 8'hfe;
      17'd73358: data = 8'hfe;
      17'd73359: data = 8'hfe;
      17'd73360: data = 8'hfe;
      17'd73361: data = 8'h00;
      17'd73362: data = 8'h00;
      17'd73363: data = 8'h00;
      17'd73364: data = 8'h00;
      17'd73365: data = 8'h00;
      17'd73366: data = 8'hfe;
      17'd73367: data = 8'h00;
      17'd73368: data = 8'hfe;
      17'd73369: data = 8'hfd;
      17'd73370: data = 8'hfe;
      17'd73371: data = 8'hfe;
      17'd73372: data = 8'h00;
      17'd73373: data = 8'hfe;
      17'd73374: data = 8'h00;
      17'd73375: data = 8'h02;
      17'd73376: data = 8'h00;
      17'd73377: data = 8'h00;
      17'd73378: data = 8'h01;
      17'd73379: data = 8'h01;
      17'd73380: data = 8'h01;
      17'd73381: data = 8'h01;
      17'd73382: data = 8'h01;
      17'd73383: data = 8'h01;
      17'd73384: data = 8'h00;
      17'd73385: data = 8'h00;
      17'd73386: data = 8'h00;
      17'd73387: data = 8'hfd;
      17'd73388: data = 8'h00;
      17'd73389: data = 8'h01;
      17'd73390: data = 8'h00;
      17'd73391: data = 8'h00;
      17'd73392: data = 8'h01;
      17'd73393: data = 8'hfe;
      17'd73394: data = 8'h00;
      17'd73395: data = 8'h00;
      17'd73396: data = 8'hfe;
      17'd73397: data = 8'hfe;
      17'd73398: data = 8'h00;
      17'd73399: data = 8'h00;
      17'd73400: data = 8'h00;
      17'd73401: data = 8'h00;
      17'd73402: data = 8'hfe;
      17'd73403: data = 8'hfe;
      17'd73404: data = 8'hfe;
      17'd73405: data = 8'hfe;
      17'd73406: data = 8'h00;
      17'd73407: data = 8'hfe;
      17'd73408: data = 8'h01;
      17'd73409: data = 8'h00;
      17'd73410: data = 8'h00;
      17'd73411: data = 8'h01;
      17'd73412: data = 8'h01;
      17'd73413: data = 8'h00;
      17'd73414: data = 8'h00;
      17'd73415: data = 8'h01;
      17'd73416: data = 8'h00;
      17'd73417: data = 8'h00;
      17'd73418: data = 8'h01;
      17'd73419: data = 8'h01;
      17'd73420: data = 8'h00;
      17'd73421: data = 8'h00;
      17'd73422: data = 8'h02;
      17'd73423: data = 8'h01;
      17'd73424: data = 8'h01;
      17'd73425: data = 8'h01;
      17'd73426: data = 8'h01;
      17'd73427: data = 8'h01;
      17'd73428: data = 8'h02;
      17'd73429: data = 8'h02;
      17'd73430: data = 8'h01;
      17'd73431: data = 8'h00;
      17'd73432: data = 8'h01;
      17'd73433: data = 8'h00;
      17'd73434: data = 8'h01;
      17'd73435: data = 8'h00;
      17'd73436: data = 8'hfe;
      17'd73437: data = 8'h01;
      17'd73438: data = 8'h00;
      17'd73439: data = 8'hfe;
      17'd73440: data = 8'h00;
      17'd73441: data = 8'h00;
      17'd73442: data = 8'h00;
      17'd73443: data = 8'h00;
      17'd73444: data = 8'hfd;
      17'd73445: data = 8'hfe;
      17'd73446: data = 8'h00;
      17'd73447: data = 8'hfd;
      17'd73448: data = 8'hfe;
      17'd73449: data = 8'hfe;
      17'd73450: data = 8'hfe;
      17'd73451: data = 8'hfd;
      17'd73452: data = 8'hfc;
      17'd73453: data = 8'hfe;
      17'd73454: data = 8'hfd;
      17'd73455: data = 8'hfe;
      17'd73456: data = 8'hfe;
      17'd73457: data = 8'hfe;
      17'd73458: data = 8'h00;
      17'd73459: data = 8'h01;
      17'd73460: data = 8'hfd;
      17'd73461: data = 8'hfe;
      17'd73462: data = 8'h00;
      17'd73463: data = 8'hfd;
      17'd73464: data = 8'hfd;
      17'd73465: data = 8'hfe;
      17'd73466: data = 8'hfd;
      17'd73467: data = 8'h00;
      17'd73468: data = 8'h01;
      17'd73469: data = 8'hfe;
      17'd73470: data = 8'h00;
      17'd73471: data = 8'h02;
      17'd73472: data = 8'h01;
      17'd73473: data = 8'h01;
      17'd73474: data = 8'h01;
      17'd73475: data = 8'hfe;
      17'd73476: data = 8'h00;
      17'd73477: data = 8'hfe;
      17'd73478: data = 8'hfd;
      17'd73479: data = 8'hfe;
      17'd73480: data = 8'hfd;
      17'd73481: data = 8'hfc;
      17'd73482: data = 8'hfd;
      17'd73483: data = 8'hfe;
      17'd73484: data = 8'hfd;
      17'd73485: data = 8'h00;
      17'd73486: data = 8'h01;
      17'd73487: data = 8'h00;
      17'd73488: data = 8'h00;
      17'd73489: data = 8'hfe;
      17'd73490: data = 8'hfe;
      17'd73491: data = 8'hfe;
      17'd73492: data = 8'h00;
      17'd73493: data = 8'h00;
      17'd73494: data = 8'hfd;
      17'd73495: data = 8'h01;
      17'd73496: data = 8'h01;
      17'd73497: data = 8'hfe;
      17'd73498: data = 8'h01;
      17'd73499: data = 8'h01;
      17'd73500: data = 8'h00;
      17'd73501: data = 8'h00;
      17'd73502: data = 8'h00;
      17'd73503: data = 8'h00;
      17'd73504: data = 8'hfe;
      17'd73505: data = 8'hfe;
      17'd73506: data = 8'hfe;
      17'd73507: data = 8'hfd;
      17'd73508: data = 8'hfd;
      17'd73509: data = 8'hfe;
      17'd73510: data = 8'hfe;
      17'd73511: data = 8'hfe;
      17'd73512: data = 8'hfe;
      17'd73513: data = 8'hfe;
      17'd73514: data = 8'hfd;
      17'd73515: data = 8'hfd;
      17'd73516: data = 8'hfe;
      17'd73517: data = 8'hfe;
      17'd73518: data = 8'hfe;
      17'd73519: data = 8'h00;
      17'd73520: data = 8'h00;
      17'd73521: data = 8'hfe;
      17'd73522: data = 8'hfe;
      17'd73523: data = 8'h01;
      17'd73524: data = 8'hfe;
      17'd73525: data = 8'hfe;
      17'd73526: data = 8'h00;
      17'd73527: data = 8'hfe;
      17'd73528: data = 8'h00;
      17'd73529: data = 8'h00;
      17'd73530: data = 8'hfe;
      17'd73531: data = 8'hfe;
      17'd73532: data = 8'h00;
      17'd73533: data = 8'h00;
      17'd73534: data = 8'h00;
      17'd73535: data = 8'h00;
      17'd73536: data = 8'h00;
      17'd73537: data = 8'h00;
      17'd73538: data = 8'hfe;
      17'd73539: data = 8'hfe;
      17'd73540: data = 8'hfe;
      17'd73541: data = 8'h00;
      17'd73542: data = 8'hfd;
      17'd73543: data = 8'hfe;
      17'd73544: data = 8'h00;
      17'd73545: data = 8'hfe;
      17'd73546: data = 8'hfe;
      17'd73547: data = 8'hfe;
      17'd73548: data = 8'h00;
      17'd73549: data = 8'h00;
      17'd73550: data = 8'h01;
      17'd73551: data = 8'hfe;
      17'd73552: data = 8'hfc;
      17'd73553: data = 8'hfe;
      17'd73554: data = 8'hfe;
      17'd73555: data = 8'hfe;
      17'd73556: data = 8'hfd;
      17'd73557: data = 8'hfd;
      17'd73558: data = 8'hfd;
      17'd73559: data = 8'hfe;
      17'd73560: data = 8'hfe;
      17'd73561: data = 8'hfe;
      17'd73562: data = 8'h01;
      17'd73563: data = 8'h02;
      17'd73564: data = 8'h01;
      17'd73565: data = 8'h01;
      17'd73566: data = 8'h01;
      17'd73567: data = 8'h00;
      17'd73568: data = 8'h00;
      17'd73569: data = 8'hfe;
      17'd73570: data = 8'hfe;
      17'd73571: data = 8'h00;
      17'd73572: data = 8'hfe;
      17'd73573: data = 8'hfe;
      17'd73574: data = 8'hfd;
      17'd73575: data = 8'hfe;
      17'd73576: data = 8'hfe;
      17'd73577: data = 8'hfe;
      17'd73578: data = 8'h00;
      17'd73579: data = 8'hfd;
      17'd73580: data = 8'hfd;
      17'd73581: data = 8'hfd;
      17'd73582: data = 8'hfc;
      17'd73583: data = 8'hfc;
      17'd73584: data = 8'hfd;
      17'd73585: data = 8'hfd;
      17'd73586: data = 8'hfd;
      17'd73587: data = 8'hfe;
      17'd73588: data = 8'hfe;
      17'd73589: data = 8'hfd;
      17'd73590: data = 8'hfd;
      17'd73591: data = 8'hfd;
      17'd73592: data = 8'hfe;
      17'd73593: data = 8'hfd;
      17'd73594: data = 8'hfd;
      17'd73595: data = 8'hfd;
      17'd73596: data = 8'hfe;
      17'd73597: data = 8'hfd;
      17'd73598: data = 8'hfd;
      17'd73599: data = 8'hfe;
      17'd73600: data = 8'hfe;
      17'd73601: data = 8'h00;
      17'd73602: data = 8'hfe;
      17'd73603: data = 8'h00;
      17'd73604: data = 8'hfe;
      17'd73605: data = 8'hfe;
      17'd73606: data = 8'hfe;
      17'd73607: data = 8'hfe;
      17'd73608: data = 8'h00;
      17'd73609: data = 8'hfe;
      17'd73610: data = 8'hfe;
      17'd73611: data = 8'h00;
      17'd73612: data = 8'h02;
      17'd73613: data = 8'h01;
      17'd73614: data = 8'h04;
      17'd73615: data = 8'h02;
      17'd73616: data = 8'h01;
      17'd73617: data = 8'h01;
      17'd73618: data = 8'h01;
      17'd73619: data = 8'h00;
      17'd73620: data = 8'hfe;
      17'd73621: data = 8'hfe;
      17'd73622: data = 8'hfe;
      17'd73623: data = 8'h01;
      17'd73624: data = 8'h00;
      17'd73625: data = 8'h01;
      17'd73626: data = 8'h01;
      17'd73627: data = 8'h02;
      17'd73628: data = 8'h01;
      17'd73629: data = 8'h01;
      17'd73630: data = 8'h02;
      17'd73631: data = 8'h01;
      17'd73632: data = 8'h00;
      17'd73633: data = 8'hfe;
      17'd73634: data = 8'hfe;
      17'd73635: data = 8'hfe;
      17'd73636: data = 8'hfe;
      17'd73637: data = 8'hfd;
      17'd73638: data = 8'hfe;
      17'd73639: data = 8'hfe;
      17'd73640: data = 8'h00;
      17'd73641: data = 8'h01;
      17'd73642: data = 8'h00;
      17'd73643: data = 8'hfe;
      17'd73644: data = 8'h00;
      17'd73645: data = 8'h00;
      17'd73646: data = 8'hfd;
      17'd73647: data = 8'hfd;
      17'd73648: data = 8'hfd;
      17'd73649: data = 8'hfa;
      17'd73650: data = 8'hfc;
      17'd73651: data = 8'hfd;
      17'd73652: data = 8'hfc;
      17'd73653: data = 8'hfd;
      17'd73654: data = 8'h00;
      17'd73655: data = 8'hfd;
      17'd73656: data = 8'hfd;
      17'd73657: data = 8'h01;
      17'd73658: data = 8'h01;
      17'd73659: data = 8'h01;
      17'd73660: data = 8'h01;
      17'd73661: data = 8'h01;
      17'd73662: data = 8'h00;
      17'd73663: data = 8'h00;
      17'd73664: data = 8'h00;
      17'd73665: data = 8'h00;
      17'd73666: data = 8'h00;
      17'd73667: data = 8'h01;
      17'd73668: data = 8'h01;
      17'd73669: data = 8'h02;
      17'd73670: data = 8'h00;
      17'd73671: data = 8'h00;
      17'd73672: data = 8'h01;
      17'd73673: data = 8'h00;
      17'd73674: data = 8'h00;
      17'd73675: data = 8'h01;
      17'd73676: data = 8'h01;
      17'd73677: data = 8'h00;
      17'd73678: data = 8'h01;
      17'd73679: data = 8'h01;
      17'd73680: data = 8'h00;
      17'd73681: data = 8'h00;
      17'd73682: data = 8'h00;
      17'd73683: data = 8'hfe;
      17'd73684: data = 8'h01;
      17'd73685: data = 8'h00;
      17'd73686: data = 8'hfe;
      17'd73687: data = 8'h01;
      17'd73688: data = 8'h01;
      17'd73689: data = 8'hfe;
      17'd73690: data = 8'h01;
      17'd73691: data = 8'h01;
      17'd73692: data = 8'hfe;
      17'd73693: data = 8'h00;
      17'd73694: data = 8'h01;
      17'd73695: data = 8'h00;
      17'd73696: data = 8'h01;
      17'd73697: data = 8'h02;
      17'd73698: data = 8'h00;
      17'd73699: data = 8'hfe;
      17'd73700: data = 8'h00;
      17'd73701: data = 8'h00;
      17'd73702: data = 8'hfe;
      17'd73703: data = 8'h01;
      17'd73704: data = 8'h00;
      17'd73705: data = 8'hfe;
      17'd73706: data = 8'h00;
      17'd73707: data = 8'hfe;
      17'd73708: data = 8'hfe;
      17'd73709: data = 8'hfe;
      17'd73710: data = 8'hfc;
      17'd73711: data = 8'hfc;
      17'd73712: data = 8'hfd;
      17'd73713: data = 8'hfa;
      17'd73714: data = 8'hfc;
      17'd73715: data = 8'hfd;
      17'd73716: data = 8'hfe;
      17'd73717: data = 8'h00;
      17'd73718: data = 8'h01;
      17'd73719: data = 8'h00;
      17'd73720: data = 8'h00;
      17'd73721: data = 8'h00;
      17'd73722: data = 8'hfe;
      17'd73723: data = 8'hfe;
      17'd73724: data = 8'hfe;
      17'd73725: data = 8'hfe;
      17'd73726: data = 8'hfe;
      17'd73727: data = 8'hfd;
      17'd73728: data = 8'hfd;
      17'd73729: data = 8'hfd;
      17'd73730: data = 8'h00;
      17'd73731: data = 8'h00;
      17'd73732: data = 8'h00;
      17'd73733: data = 8'h02;
      17'd73734: data = 8'h02;
      17'd73735: data = 8'h04;
      17'd73736: data = 8'h02;
      17'd73737: data = 8'h01;
      17'd73738: data = 8'h02;
      17'd73739: data = 8'h01;
      17'd73740: data = 8'hfe;
      17'd73741: data = 8'h00;
      17'd73742: data = 8'h01;
      17'd73743: data = 8'h01;
      17'd73744: data = 8'h01;
      17'd73745: data = 8'h02;
      17'd73746: data = 8'h01;
      17'd73747: data = 8'h02;
      17'd73748: data = 8'h04;
      17'd73749: data = 8'h01;
      17'd73750: data = 8'h01;
      17'd73751: data = 8'h01;
      17'd73752: data = 8'h00;
      17'd73753: data = 8'hfe;
      17'd73754: data = 8'hfe;
      17'd73755: data = 8'hfe;
      17'd73756: data = 8'hfd;
      17'd73757: data = 8'hfc;
      17'd73758: data = 8'hfd;
      17'd73759: data = 8'hfc;
      17'd73760: data = 8'hfe;
      17'd73761: data = 8'h00;
      17'd73762: data = 8'h00;
      17'd73763: data = 8'hfe;
      17'd73764: data = 8'h00;
      17'd73765: data = 8'hfe;
      17'd73766: data = 8'hfe;
      17'd73767: data = 8'hfe;
      17'd73768: data = 8'hfe;
      17'd73769: data = 8'hfe;
      17'd73770: data = 8'hfe;
      17'd73771: data = 8'hfd;
      17'd73772: data = 8'hfe;
      17'd73773: data = 8'hfe;
      17'd73774: data = 8'hfd;
      17'd73775: data = 8'hfe;
      17'd73776: data = 8'hfe;
      17'd73777: data = 8'h00;
      17'd73778: data = 8'hfe;
      17'd73779: data = 8'h00;
      17'd73780: data = 8'h00;
      17'd73781: data = 8'h01;
      17'd73782: data = 8'h02;
      17'd73783: data = 8'h00;
      17'd73784: data = 8'h01;
      17'd73785: data = 8'h02;
      17'd73786: data = 8'h01;
      17'd73787: data = 8'h00;
      17'd73788: data = 8'h00;
      17'd73789: data = 8'hfe;
      17'd73790: data = 8'hfe;
      17'd73791: data = 8'h00;
      17'd73792: data = 8'h00;
      17'd73793: data = 8'hfe;
      17'd73794: data = 8'h00;
      17'd73795: data = 8'h00;
      17'd73796: data = 8'h00;
      17'd73797: data = 8'h00;
      17'd73798: data = 8'h00;
      17'd73799: data = 8'h00;
      17'd73800: data = 8'hfe;
      17'd73801: data = 8'hfe;
      17'd73802: data = 8'hfd;
      17'd73803: data = 8'hfe;
      17'd73804: data = 8'hfd;
      17'd73805: data = 8'hfd;
      17'd73806: data = 8'hfd;
      17'd73807: data = 8'hfc;
      17'd73808: data = 8'hfd;
      17'd73809: data = 8'hfe;
      17'd73810: data = 8'hfd;
      17'd73811: data = 8'hfd;
      17'd73812: data = 8'hfd;
      17'd73813: data = 8'hfe;
      17'd73814: data = 8'hfd;
      17'd73815: data = 8'hfd;
      17'd73816: data = 8'hfe;
      17'd73817: data = 8'hfd;
      17'd73818: data = 8'hfd;
      17'd73819: data = 8'hfe;
      17'd73820: data = 8'hfd;
      17'd73821: data = 8'hfd;
      17'd73822: data = 8'h00;
      17'd73823: data = 8'hfe;
      17'd73824: data = 8'hfe;
      17'd73825: data = 8'hfe;
      17'd73826: data = 8'hfd;
      17'd73827: data = 8'hfe;
      17'd73828: data = 8'hfe;
      17'd73829: data = 8'h00;
      17'd73830: data = 8'h00;
      17'd73831: data = 8'h00;
      17'd73832: data = 8'h00;
      17'd73833: data = 8'hfe;
      17'd73834: data = 8'hfe;
      17'd73835: data = 8'hfe;
      17'd73836: data = 8'hfd;
      17'd73837: data = 8'hfd;
      17'd73838: data = 8'hfd;
      17'd73839: data = 8'hfc;
      17'd73840: data = 8'hfd;
      17'd73841: data = 8'hfd;
      17'd73842: data = 8'hfe;
      17'd73843: data = 8'h00;
      17'd73844: data = 8'hfe;
      17'd73845: data = 8'hfe;
      17'd73846: data = 8'hfe;
      17'd73847: data = 8'hfe;
      17'd73848: data = 8'hfe;
      17'd73849: data = 8'hfe;
      17'd73850: data = 8'hfe;
      17'd73851: data = 8'hfe;
      17'd73852: data = 8'hfe;
      17'd73853: data = 8'hfd;
      17'd73854: data = 8'hfd;
      17'd73855: data = 8'h00;
      17'd73856: data = 8'h00;
      17'd73857: data = 8'h00;
      17'd73858: data = 8'h01;
      17'd73859: data = 8'h02;
      17'd73860: data = 8'h01;
      17'd73861: data = 8'h01;
      17'd73862: data = 8'h01;
      17'd73863: data = 8'h00;
      17'd73864: data = 8'h00;
      17'd73865: data = 8'hfe;
      17'd73866: data = 8'h00;
      17'd73867: data = 8'h00;
      17'd73868: data = 8'h01;
      17'd73869: data = 8'h00;
      17'd73870: data = 8'h00;
      17'd73871: data = 8'hfe;
      17'd73872: data = 8'hfe;
      17'd73873: data = 8'h00;
      17'd73874: data = 8'h00;
      17'd73875: data = 8'h00;
      17'd73876: data = 8'hfe;
      17'd73877: data = 8'h00;
      17'd73878: data = 8'h00;
      17'd73879: data = 8'h00;
      17'd73880: data = 8'h01;
      17'd73881: data = 8'hfe;
      17'd73882: data = 8'hfd;
      17'd73883: data = 8'hfe;
      17'd73884: data = 8'hfe;
      17'd73885: data = 8'h00;
      17'd73886: data = 8'h00;
      17'd73887: data = 8'h00;
      17'd73888: data = 8'h01;
      17'd73889: data = 8'h01;
      17'd73890: data = 8'hfe;
      17'd73891: data = 8'hfe;
      17'd73892: data = 8'hfe;
      17'd73893: data = 8'hfe;
      17'd73894: data = 8'hfd;
      17'd73895: data = 8'hfd;
      17'd73896: data = 8'hfe;
      17'd73897: data = 8'hfd;
      17'd73898: data = 8'hfc;
      17'd73899: data = 8'hfe;
      17'd73900: data = 8'hfe;
      17'd73901: data = 8'hfd;
      17'd73902: data = 8'hfe;
      17'd73903: data = 8'hfd;
      17'd73904: data = 8'hfe;
      17'd73905: data = 8'h00;
      17'd73906: data = 8'hfe;
      17'd73907: data = 8'hfe;
      17'd73908: data = 8'hfe;
      17'd73909: data = 8'hfe;
      17'd73910: data = 8'hfd;
      17'd73911: data = 8'hfd;
      17'd73912: data = 8'hfe;
      17'd73913: data = 8'hfd;
      17'd73914: data = 8'hfe;
      17'd73915: data = 8'hfe;
      17'd73916: data = 8'h00;
      17'd73917: data = 8'h00;
      17'd73918: data = 8'h00;
      17'd73919: data = 8'h01;
      17'd73920: data = 8'h01;
      17'd73921: data = 8'h00;
      17'd73922: data = 8'h00;
      17'd73923: data = 8'h00;
      17'd73924: data = 8'h00;
      17'd73925: data = 8'hfe;
      17'd73926: data = 8'h00;
      17'd73927: data = 8'hfe;
      17'd73928: data = 8'hfe;
      17'd73929: data = 8'h00;
      17'd73930: data = 8'h01;
      17'd73931: data = 8'h02;
      17'd73932: data = 8'h02;
      17'd73933: data = 8'h02;
      17'd73934: data = 8'h01;
      17'd73935: data = 8'h02;
      17'd73936: data = 8'h00;
      17'd73937: data = 8'h00;
      17'd73938: data = 8'hfd;
      17'd73939: data = 8'hfd;
      17'd73940: data = 8'hfe;
      17'd73941: data = 8'hfd;
      17'd73942: data = 8'hfe;
      17'd73943: data = 8'hfe;
      17'd73944: data = 8'hfe;
      17'd73945: data = 8'hfe;
      17'd73946: data = 8'hfd;
      17'd73947: data = 8'h00;
      17'd73948: data = 8'hfe;
      17'd73949: data = 8'h00;
      17'd73950: data = 8'hfe;
      17'd73951: data = 8'h00;
      17'd73952: data = 8'h00;
      17'd73953: data = 8'h00;
      17'd73954: data = 8'h00;
      17'd73955: data = 8'hfe;
      17'd73956: data = 8'h00;
      17'd73957: data = 8'hfe;
      17'd73958: data = 8'hfe;
      17'd73959: data = 8'h00;
      17'd73960: data = 8'h00;
      17'd73961: data = 8'h02;
      17'd73962: data = 8'h01;
      17'd73963: data = 8'h02;
      17'd73964: data = 8'h01;
      17'd73965: data = 8'h01;
      17'd73966: data = 8'h01;
      17'd73967: data = 8'h00;
      17'd73968: data = 8'h01;
      17'd73969: data = 8'h01;
      17'd73970: data = 8'h00;
      17'd73971: data = 8'h01;
      17'd73972: data = 8'h01;
      17'd73973: data = 8'h00;
      17'd73974: data = 8'h00;
      17'd73975: data = 8'h02;
      17'd73976: data = 8'h01;
      17'd73977: data = 8'h00;
      17'd73978: data = 8'h01;
      17'd73979: data = 8'h01;
      17'd73980: data = 8'h01;
      17'd73981: data = 8'h01;
      17'd73982: data = 8'h01;
      17'd73983: data = 8'h01;
      17'd73984: data = 8'h00;
      17'd73985: data = 8'h00;
      17'd73986: data = 8'h00;
      17'd73987: data = 8'hfe;
      17'd73988: data = 8'h00;
      17'd73989: data = 8'h00;
      17'd73990: data = 8'h00;
      17'd73991: data = 8'h00;
      17'd73992: data = 8'h01;
      17'd73993: data = 8'h00;
      17'd73994: data = 8'hfe;
      17'd73995: data = 8'h00;
      17'd73996: data = 8'h02;
      17'd73997: data = 8'hfe;
      17'd73998: data = 8'hfe;
      17'd73999: data = 8'h00;
      17'd74000: data = 8'hfe;
      17'd74001: data = 8'hfe;
      17'd74002: data = 8'hfe;
      17'd74003: data = 8'hfe;
      17'd74004: data = 8'hfd;
      17'd74005: data = 8'hfe;
      17'd74006: data = 8'hfe;
      17'd74007: data = 8'h00;
      17'd74008: data = 8'hfe;
      17'd74009: data = 8'hfe;
      17'd74010: data = 8'hfd;
      17'd74011: data = 8'hfd;
      17'd74012: data = 8'hfd;
      17'd74013: data = 8'hfd;
      17'd74014: data = 8'hfd;
      17'd74015: data = 8'hfd;
      17'd74016: data = 8'hfd;
      17'd74017: data = 8'hfd;
      17'd74018: data = 8'hfe;
      17'd74019: data = 8'hfe;
      17'd74020: data = 8'h00;
      17'd74021: data = 8'h00;
      17'd74022: data = 8'h00;
      17'd74023: data = 8'h01;
      17'd74024: data = 8'h01;
      17'd74025: data = 8'hfe;
      17'd74026: data = 8'hfe;
      17'd74027: data = 8'hfd;
      17'd74028: data = 8'hfe;
      17'd74029: data = 8'h00;
      17'd74030: data = 8'h00;
      17'd74031: data = 8'hfe;
      17'd74032: data = 8'h00;
      17'd74033: data = 8'h01;
      17'd74034: data = 8'h00;
      17'd74035: data = 8'hfe;
      17'd74036: data = 8'h00;
      17'd74037: data = 8'h00;
      17'd74038: data = 8'h00;
      17'd74039: data = 8'h00;
      17'd74040: data = 8'hfd;
      17'd74041: data = 8'hfd;
      17'd74042: data = 8'hfe;
      17'd74043: data = 8'hfd;
      17'd74044: data = 8'hfe;
      17'd74045: data = 8'hfe;
      17'd74046: data = 8'hfe;
      17'd74047: data = 8'hfe;
      17'd74048: data = 8'h00;
      17'd74049: data = 8'h00;
      17'd74050: data = 8'h00;
      17'd74051: data = 8'h00;
      17'd74052: data = 8'h00;
      17'd74053: data = 8'h00;
      17'd74054: data = 8'h01;
      17'd74055: data = 8'hfe;
      17'd74056: data = 8'hfe;
      17'd74057: data = 8'hfe;
      17'd74058: data = 8'hfc;
      17'd74059: data = 8'hfd;
      17'd74060: data = 8'h00;
      17'd74061: data = 8'hfe;
      17'd74062: data = 8'hfe;
      17'd74063: data = 8'h00;
      17'd74064: data = 8'h00;
      17'd74065: data = 8'h00;
      17'd74066: data = 8'h00;
      17'd74067: data = 8'h01;
      17'd74068: data = 8'h00;
      17'd74069: data = 8'hfe;
      17'd74070: data = 8'hfc;
      17'd74071: data = 8'hfc;
      17'd74072: data = 8'hfc;
      17'd74073: data = 8'hfa;
      17'd74074: data = 8'hfa;
      17'd74075: data = 8'hfc;
      17'd74076: data = 8'hfd;
      17'd74077: data = 8'hfe;
      17'd74078: data = 8'h00;
      17'd74079: data = 8'h00;
      17'd74080: data = 8'h01;
      17'd74081: data = 8'h01;
      17'd74082: data = 8'h01;
      17'd74083: data = 8'h01;
      17'd74084: data = 8'h00;
      17'd74085: data = 8'h00;
      17'd74086: data = 8'h00;
      17'd74087: data = 8'hfe;
      17'd74088: data = 8'h00;
      17'd74089: data = 8'hfe;
      17'd74090: data = 8'hfd;
      17'd74091: data = 8'h00;
      17'd74092: data = 8'h00;
      17'd74093: data = 8'h01;
      17'd74094: data = 8'h02;
      17'd74095: data = 8'h02;
      17'd74096: data = 8'h02;
      17'd74097: data = 8'h04;
      17'd74098: data = 8'h02;
      17'd74099: data = 8'h00;
      17'd74100: data = 8'h00;
      17'd74101: data = 8'h00;
      17'd74102: data = 8'h01;
      17'd74103: data = 8'h00;
      17'd74104: data = 8'hfe;
      17'd74105: data = 8'hfe;
      17'd74106: data = 8'h00;
      17'd74107: data = 8'h01;
      17'd74108: data = 8'h01;
      17'd74109: data = 8'h01;
      17'd74110: data = 8'h01;
      17'd74111: data = 8'h02;
      17'd74112: data = 8'h00;
      17'd74113: data = 8'h00;
      17'd74114: data = 8'h00;
      17'd74115: data = 8'h00;
      17'd74116: data = 8'hfe;
      17'd74117: data = 8'hfd;
      17'd74118: data = 8'hfd;
      17'd74119: data = 8'hfd;
      17'd74120: data = 8'hfd;
      17'd74121: data = 8'hfe;
      17'd74122: data = 8'h01;
      17'd74123: data = 8'h01;
      17'd74124: data = 8'h04;
      17'd74125: data = 8'h02;
      17'd74126: data = 8'h02;
      17'd74127: data = 8'h02;
      17'd74128: data = 8'h02;
      17'd74129: data = 8'h00;
      17'd74130: data = 8'h00;
      17'd74131: data = 8'h00;
      17'd74132: data = 8'hfe;
      17'd74133: data = 8'h01;
      17'd74134: data = 8'h01;
      17'd74135: data = 8'h00;
      17'd74136: data = 8'h01;
      17'd74137: data = 8'h00;
      17'd74138: data = 8'h01;
      17'd74139: data = 8'h01;
      17'd74140: data = 8'h01;
      17'd74141: data = 8'h00;
      17'd74142: data = 8'hfe;
      17'd74143: data = 8'h00;
      17'd74144: data = 8'h00;
      17'd74145: data = 8'h00;
      17'd74146: data = 8'hfe;
      17'd74147: data = 8'hfe;
      17'd74148: data = 8'h00;
      17'd74149: data = 8'hfe;
      17'd74150: data = 8'hfe;
      17'd74151: data = 8'h00;
      17'd74152: data = 8'h01;
      17'd74153: data = 8'h00;
      17'd74154: data = 8'h00;
      17'd74155: data = 8'h01;
      17'd74156: data = 8'h01;
      17'd74157: data = 8'hfe;
      17'd74158: data = 8'h00;
      17'd74159: data = 8'h00;
      17'd74160: data = 8'hfe;
      17'd74161: data = 8'h00;
    endcase
  end
endmodule
